// Created by: vgen.pl 
module vgen (clk, check, done);
   input clk;
   input check;
   output done;
   initial $write("\n*** Vgen.v starting, seed = 5\n");
   // verilator lint_off UNSIGNED
   // verilator lint_off CMPCONST
   // verilator lint_off WIDTH

   reg signed [127:  0] W0001                     ; //=128'hffffffffffffffffffffffffffffffff
   reg        [  3:  0] W0002                     ; //=4'h0
   reg signed [127:  0] W0003 /*verilator public*/; //=128'hffffffffffffffffffffffffffffffff
   reg        [118:  0] W0004 /*verilator public*/; //=119'h2f54d600000000ffffffff00000000
   reg        [  2:  0] W0005 /*verilator public*/; //=3'h1
   reg signed [ 35:  0] W0006 /*verilator public*/; //=36'h000000001
   reg signed [ 94:  0] W0007                     ; //=95'h1feb10faffffffff00000000
   reg        [ 60:  0] W0008 /*verilator public*/; //=61'h1fffffffffffffff
   reg signed [101:  0] W0009 /*verilator public*/; //=102'h00000000000000000000000000
   reg signed [ 62:  0] W0010                     ; //=63'h0000000000000001
   reg        [  6:  0] W0011                     ; //=7'h7f
   reg        [108:  0] W0012 /*verilator public*/; //=109'h1fffffffffffffffffffffffffff
   reg        [108:  0] W0013                     ; //=109'h1fffffffffffffffffffffffffff
   reg        [ 66:  0] W0014                     ; //=67'h00000000000000000
   reg signed [  7:  0] W0015                     ; //=8'h00
   reg signed [ 87:  0] W0016 /*verilator public*/; //=88'h0000000000000000000000
   reg signed [ 31:  0] W0017 /*verilator public*/; //=32'hffffffff
   reg signed [123:  0] W0018                     ; //=124'h0000000000000000000000000000000
   reg signed [ 96:  0] W0019                     ; //=97'h000000001abf37a3000000001
   reg signed [ 96:  0] W0020                     ; //=97'h1ffffffffffffffffffffffff
   reg signed [125:  0] W0021 /*verilator public*/; //=126'h3fffffffffffffffffffffffffffffff
   reg signed [122:  0] W0022                     ; //=123'h7ffffffbce03e2bdb14609fe7e28b41
   reg signed [ 83:  0] W0023                     ; //=84'h0000000000000e1fe9094
   reg signed [ 83:  0] W0024                     ; //=84'h0f66afffffffe308b3d7c
   reg        [ 74:  0] W0025                     ; //=75'h0000000000000000000
   reg signed [ 38:  0] W0026                     ; //=39'h005f38482c
   reg signed [  6:  0] W0027                     ; //=7'h7f
   reg signed [ 38:  0] W0028                     ; //=39'h005f38482c
   reg signed [ 94:  0] W0029                     ; //=95'h000000000000000000000000
   reg signed [ 94:  0] W0030                     ; //=95'h3691dbd700000000ffffffff
   reg signed [ 63:  0] W0031                     ; //=64'hfffffffe00000001
   reg signed [ 63:  0] W0032                     ; //=64'hfffffffe00000001
   reg        [ 31:  0] W0033 /*verilator public*/; //=32'hffffffff
   reg        [ 94:  0] W0034 /*verilator public*/; //=95'h7fffffffdccdbaa8bfb519ef
   reg signed [ 89:  0] W0035 /*verilator public*/; //=90'h0000000ae9a2f0b00000000
   reg        [ 94:  0] W0036                     ; //=95'h7fffffffdccdbaa8bfb519ef
   reg signed [ 30:  0] W0037                     ; //=31'h7fffffff
   reg signed [  2:  0] W0038                     ; //=3'h0
   reg signed [ 66:  0] W0039                     ; //=67'h200000001fc7de7a7
   reg signed [  3:  0] W0040                     ; //=4'h0
   reg signed [ 30:  0] W0041                     ; //=31'h00000000
   reg signed [  6:  0] W0042                     ; //=7'h7f
   reg signed [ 98:  0] W0043                     ; //=99'h7ffffffffffffffffffffffff
   reg        [ 84:  0] W0044                     ; //=85'h0000000000000000000000
   reg        [106:  0] W0045                     ; //=107'h000000000000000000000000000
   reg        [ 84:  0] W0046                     ; //=85'h0000000000000000000000
   reg signed [ 95:  0] W0047                     ; //=96'hffffffffffffffffffffffff
   reg        [ 62:  0] W0048                     ; //=63'h00000001bf003b47
   reg signed [ 50:  0] W0049                     ; //=51'h0000000000000
   reg signed [107:  0] W0050                     ; //=108'h0170f5f330fffffffff5d6adc0b
   reg signed [107:  0] W0051                     ; //=108'h0170f5f330fffffffff5d6adc0b
   reg signed [  1:  0] W0052 /*verilator public*/; //=2'h0
   reg signed [  1:  0] W0053                     ; //=2'h0
   reg signed [  1:  0] W0054 /*verilator public*/; //=2'h0
   reg signed [ 70:  0] W0055                     ; //=71'h000000000000000000
   reg signed [ 19:  0] W0056                     ; //=20'h00000
   reg        [ 52:  0] W0057                     ; //=53'h0a9dcf00000001
   reg        [ 98:  0] W0058                     ; //=99'h0000000000000000000000000
   reg signed [ 84:  0] W0059                     ; //=85'h1fffffffffffffc422fb6e
   reg        [127:  0] W0060                     ; //=128'h00000000000000000000000000000000
   reg        [  0:  0] W0061                     ; //=1'h1
   reg signed [ 60:  0] W0062                     ; //=61'h1fffffffffffffff
   reg signed [ 27:  0] W0063                     ; //=28'h0000000
   reg signed [ 24:  0] W0064                     ; //=25'h1ffffff
   reg signed [127:  0] W0065                     ; //=128'hffffffffffffffffffffffffffffffff
   reg signed [  7:  0] W0066                     ; //=8'h00
   reg        [ 50:  0] W0067                     ; //=51'h0000000000000
   reg signed [ 14:  0] W0068                     ; //=15'h0000
   reg        [122:  0] W0069 /*verilator public*/; //=123'h0000000000000000000000000000000
   reg        [122:  0] W0070                     ; //=123'h0000000000000000000000000000000
   reg        [122:  0] W0071                     ; //=123'h0000000000000000000000000000000
   reg signed [125:  0] W0072                     ; //=126'h00000000000000000000000000000000
   reg signed [ 50:  0] W0073                     ; //=51'h7ffffffffffff
   reg signed [ 38:  0] W0074                     ; //=39'h0000000000
   reg        [125:  0] W0075                     ; //=126'h00000000000000000000000000000000
   reg        [125:  0] W0076                     ; //=126'h00000000000000000000000000000000
   reg signed [ 98:  0] W0077                     ; //=99'h7ffffffffffffffffffffffff
   reg        [ 23:  0] W0078                     ; //=24'hffffff
   reg        [125:  0] W0079                     ; //=126'h00000000000000000000000000000000
   reg        [  7:  0] W0080                     ; //=8'h00
   reg signed [110:  0] W0081 /*verilator public*/; //=111'h5d8cffffffff9b20638fffffffff
   reg signed [ 13:  0] W0082 /*verilator public*/; //=14'h0000
   reg signed [ 31:  0] W0083                     ; //=32'h00000000
   reg signed [  5:  0] W0084                     ; //=6'h30
   reg signed [ 89:  0] W0085 /*verilator public*/; //=90'h3ffffffffffffffffffffff
   reg signed [ 50:  0] W0086                     ; //=51'h0000000000000
   reg signed [ 25:  0] W0087                     ; //=26'h0000001
   reg        [ 67:  0] W0088 /*verilator public*/; //=68'h00000000000000000
   reg signed [ 78:  0] W0089                     ; //=79'h00000000000000000000
   reg signed [  5:  0] W0090                     ; //=6'h1b
   reg signed [ 77:  0] W0091 /*verilator public*/; //=78'h3fffffffffffffffffff
   reg signed [ 77:  0] W0092                     ; //=78'h3fffffffffffffffffff
   reg signed [127:  0] W0093                     ; //=128'hffffffffffffffffffffffffffffffff
   reg signed [126:  0] W0094                     ; //=127'h00000000000000000000000000000000
   reg signed [ 18:  0] W0095                     ; //=19'h7ffff
   reg signed [  7:  0] W0096                     ; //=8'h00
   reg signed [127:  0] W0097                     ; //=128'hffffffffffffffffffffffffffffffff
   reg signed [127:  0] W0098                     ; //=128'hffffffffffffffffffffffffffffffff
   reg signed [ 19:  0] W0099 /*verilator public*/; //=20'h00000
   reg signed [ 19:  0] W0100                     ; //=20'hfffff
   reg signed [ 74:  0] W0101 /*verilator public*/; //=75'h7ff7e019ac646679f3d
   reg signed [ 85:  0] W0102                     ; //=86'h3fffffffffffffffffffff
   reg signed [121:  0] W0103                     ; //=122'h3ffffffffffffffffffffffffffffff
   reg signed [121:  0] W0104                     ; //=122'h3ffffffffffffffffffffffffffffff
   reg signed [  3:  0] W0105                     ; //=4'h0
   reg signed [ 88:  0] W0106                     ; //=89'h0000000fb47be1e00000001
   reg signed [ 88:  0] W0107 /*verilator public*/; //=89'h1ffffff04b841e1ffffffff
   reg signed [ 66:  0] W0108                     ; //=67'h00000000000000000
   reg signed [ 66:  0] W0109                     ; //=67'h00000000000000000
   reg signed [ 60:  0] W0110                     ; //=61'h0000000000000000
   reg signed [  6:  0] W0111                     ; //=7'h01
   reg        [ 39:  0] W0112                     ; //=40'h0000000000
   reg        [ 39:  0] W0113                     ; //=40'h0000000000
   reg signed [ 78:  0] W0114                     ; //=79'h0001ffffffff00000000
   reg signed [ 78:  0] W0115 /*verilator public*/; //=79'h0001ffffffff00000000
   reg        [ 80:  0] W0116                     ; //=81'h000000000000000000001
   reg signed [ 87:  0] W0117                     ; //=88'h0000000000000000000000
   reg signed [ 87:  0] W0118                     ; //=88'h0000000000000000000000
   reg        [ 98:  0] W0119                     ; //=99'h0ffffffffdc3c268800000000
   reg        [  0:  0] W0120                     ; //=1'h0
   reg        [ 39:  0] W0121                     ; //=40'h0000000000
   reg signed [ 37:  0] W0122                     ; //=38'h0000000000
   reg signed [ 45:  0] W0123                     ; //=46'h000000000000
   reg        [ 70:  0] W0124 /*verilator public*/; //=71'h7fffffffffffffffff
   reg        [  7:  0] W0125 /*verilator public*/; //=8'h00
   reg signed [ 82:  0] W0126                     ; //=83'h7ffff00000000397f927d
   reg signed [ 75:  0] W0127                     ; //=76'hfffffffffffffffffff
   reg signed [ 14:  0] W0128                     ; //=15'h0000
   reg        [ 51:  0] W0129                     ; //=52'hfffffffffffff
   reg signed [127:  0] W0130 /*verilator public*/; //=128'hffffffffffffffffffffffffffffffff
   reg signed [ 66:  0] W0131                     ; //=67'h00000000000000001
   reg signed [125:  0] W0132                     ; //=126'h3ee9a075ffffffffef0f331858d8680b
   reg signed [ 62:  0] W0133                     ; //=63'h7fffffffffffffff
   reg        [ 39:  0] W0134                     ; //=40'hffffffffff
   reg signed [111:  0] W0135                     ; //=112'hffffffffffffffffffffffffffff
   reg        [ 76:  0] W0136                     ; //=77'h00000000000000000000
   reg        [  0:  0] W0137 /*verilator public*/; //=1'h1
   reg        [113:  0] W0138                     ; //=114'h3ffffffffffffffffffffffffffff
   reg signed [114:  0] W0139                     ; //=115'h7ffffffffffffffffffffffffffff
   reg signed [ 41:  0] W0140 /*verilator public*/; //=42'h00000000000
   reg signed [  6:  0] W0141 /*verilator public*/; //=7'h7f
   reg        [126:  0] W0142                     ; //=127'h00000000000000000000000000000000
   reg signed [127:  0] W0143 /*verilator public*/; //=128'h00000000000000000000000000000000
   reg signed [ 90:  0] W0144 /*verilator public*/; //=91'h0fc147500000000a1a6dc1c
   reg signed [ 90:  0] W0145                     ; //=91'h0fc147500000000a1a6dc1c
   reg signed [ 52:  0] W0146                     ; //=53'h1fffffffffffff
   reg signed [ 75:  0] W0147                     ; //=76'hbc2ffffffff61887cef
   reg signed [ 95:  0] W0148                     ; //=96'hfffffffffffffffffffffffe
   reg signed [ 95:  0] W0149                     ; //=96'hfffffffffffffffffffffffe
   reg signed [ 94:  0] W0150                     ; //=95'h496e2428ffffffff00000001
   reg signed [  5:  0] W0151 /*verilator public*/; //=6'h00
   reg        [ 31:  0] W0152 /*verilator public*/; //=32'he0000000
   reg signed [ 34:  0] W0153                     ; //=35'h700000000
   reg signed [ 34:  0] W0154                     ; //=35'h700000000
   reg signed [ 34:  0] W0155                     ; //=35'h000000000
   reg signed [120:  0] W0156                     ; //=121'h000000003d719e8ffffffffffffffff
   reg        [106:  0] W0157                     ; //=107'h000000000000000000000000000
   reg signed [107:  0] W0158 /*verilator public*/; //=108'h000000000000000000000000001
   reg signed [ 59:  0] W0159                     ; //=60'h000000000000001
   reg        [  6:  0] W0160                     ; //=7'h7f
   reg        [ 95:  0] W0161 /*verilator public*/; //=96'hfffffffffffffffffffffffd
   reg signed [116:  0] W0162                     ; //=117'h1fffffffffffffffffffffffffffff
   reg        [ 86:  0] W0163 /*verilator public*/; //=87'h7fffffffffffffffffffff
   reg signed [127:  0] W0164 /*verilator public*/; //=128'hffffffffffffffffffffffffffffffff
   reg        [ 64:  0] W0165                     ; //=65'h00000000004000000
   reg signed [ 86:  0] W0166 /*verilator public*/; //=87'h0000000000000000000000
   reg signed [ 17:  0] W0167 /*verilator public*/; //=18'h00002
   reg signed [ 17:  0] W0168                     ; //=18'h00002
   reg signed [ 95:  0] W0169                     ; //=96'h2eb5a3fd79a326f8a74f99be
   reg signed [117:  0] W0170                     ; //=118'h3fffffffffffffffffffffffffffff
   reg signed [ 96:  0] W0171                     ; //=97'h1ffffffffffffffffffffffff
   reg        [ 94:  0] W0172 /*verilator public*/; //=95'h000000000000000000000000
   reg        [116:  0] W0173 /*verilator public*/; //=117'h000000000000000000000000000000
   reg        [116:  0] W0174                     ; //=117'h1fffffffffffffffffffffffffffff
   reg        [ 22:  0] W0175                     ; //=23'h000000
   reg        [  0:  0] W0176                     ; //=1'h1
   reg        [ 37:  0] W0177 /*verilator public*/; //=38'h3c00000003
   reg signed [ 67:  0] W0178 /*verilator public*/; //=68'hf00000000ffffffff
   reg signed [ 67:  0] W0179                     ; //=68'h00000000000000000
   reg signed [  7:  0] W0180                     ; //=8'hff
   reg        [ 34:  0] W0181                     ; //=35'h7ffffffff
   reg signed [127:  0] W0182                     ; //=128'hffffffffffffffffffffffffffffffff
   reg signed [ 58:  0] W0183                     ; //=59'h7ffffffffffffff
   reg        [ 42:  0] W0184                     ; //=43'h7ffffffffff
   reg        [  4:  0] W0185 /*verilator public*/; //=5'h01
   reg        [119:  0] W0186 /*verilator public*/; //=120'h000000000000000000000000000000
   reg signed [120:  0] W0187 /*verilator public*/; //=121'h1ffffff000000000000000064c42d4b
   reg signed [127:  0] W0188                     ; //=128'h00000000000000000000000000000000
   reg        [104:  0] W0189 /*verilator public*/; //=105'h1ffffffc1e7d361800000002660
   reg signed [122:  0] W0190                     ; //=123'h7ffffff079f4d86000000009983636f
   reg        [  8:  0] W0191                     ; //=9'h000
   reg signed [  2:  0] W0192                     ; //=3'h7
   reg signed [  1:  0] W0193                     ; //=2'h0
   reg signed [ 34:  0] W0194                     ; //=35'h600000000
   reg signed [ 30:  0] W0195                     ; //=31'h00000000
   reg        [  0:  0] W0196                     ; //=1'h1
   reg signed [110:  0] W0197                     ; //=111'h0000000000000000000000000000
   reg        [ 14:  0] W0198                     ; //=15'h0000
   reg signed [ 24:  0] W0199 /*verilator public*/; //=25'h1930f53
   reg        [  0:  0] W0200                     ; //=1'h0
   reg signed [ 61:  0] W0201 /*verilator public*/; //=62'h3fffffffffffffff
   reg signed [127:  0] W0202                     ; //=128'h00000000000000000000000000000000
   reg        [ 82:  0] W0203                     ; //=83'h7b3155312a8ed00000000
   reg        [ 28:  0] W0204                     ; //=29'h1f3fc1c3
   reg        [  3:  0] W0205                     ; //=4'h0
   reg signed [ 98:  0] W0206                     ; //=99'h0000000000000000000000000
   reg signed [124:  0] W0207                     ; //=125'h00000000000000000000000000000001
   reg signed [104:  0] W0208                     ; //=105'h000000000000000000000000000
   reg signed [100:  0] W0209                     ; //=101'h1fffffffff0000000000000001
   reg        [  1:  0] W0210                     ; //=2'h0
   reg signed [110:  0] W0211 /*verilator public*/; //=111'h0000000000000000000000000000
   reg        [ 62:  0] W0212 /*verilator public*/; //=63'h7fffffffffffffff
   reg signed [ 97:  0] W0213                     ; //=98'h0000000000000000000000001
   reg signed [100:  0] W0214 /*verilator public*/; //=101'h1fffffffff0000000000000001
   reg        [  5:  0] W0215                     ; //=6'h00
   reg        [ 14:  0] W0216 /*verilator public*/; //=15'h0000
   reg signed [102:  0] W0217                     ; //=103'h00000000000000000000000000
   reg signed [102:  0] W0218                     ; //=103'h0085bac6fde88fbe57a202d84c
   reg signed [102:  0] W0219 /*verilator public*/; //=103'h00000000000000000000000001
   reg signed [ 34:  0] W0220 /*verilator public*/; //=35'h0fffffffe
   reg signed [104:  0] W0221                     ; //=105'h18b7e03b2359874995a00000000
   reg signed [ 98:  0] W0222                     ; //=99'h0000000000000000000000000
   reg        [124:  0] W0223 /*verilator public*/; //=125'h04000000000000000000000000000000
   reg        [ 98:  0] W0224                     ; //=99'h7ffffffffffffffffffffffff
   reg signed [102:  0] W0225                     ; //=103'h7fffffffffffffffffffffffff
   reg signed [  4:  0] W0226                     ; //=5'h00
   reg signed [  4:  0] W0227                     ; //=5'h1f
   reg signed [  4:  0] W0228                     ; //=5'h10
   reg signed [  2:  0] W0229 /*verilator public*/; //=3'h3
   reg        [  0:  0] W0230                     ; //=1'h0
   reg        [127:  0] W0231                     ; //=128'h00000000000000000000000000000000
   reg        [ 94:  0] W0232                     ; //=95'h000000000000000000000000
   reg signed [ 13:  0] W0233                     ; //=14'h0000
   reg signed [126:  0] W0234 /*verilator public*/; //=127'h00000000000000000000000000000000
   reg signed [  7:  0] W0235                     ; //=8'hff
   reg signed [ 36:  0] W0236 /*verilator public*/; //=37'h1fffffffff
   reg        [  0:  0] W0237                     ; //=1'h0
   reg signed [118:  0] W0238                     ; //=119'h7fffff00000000ffffffffffffffff
   reg signed [122:  0] W0239                     ; //=123'h53fb225d8fa2187ffffffffffffffff
   reg signed [ 49:  0] W0240                     ; //=50'h0000000000000
   reg signed [ 66:  0] W0241                     ; //=67'h7ffffffffee0efff1
   reg signed [  5:  0] W0242 /*verilator public*/; //=6'h3f
   reg        [ 31:  0] W0243                     ; //=32'hffffffff
   reg signed [  7:  0] W0244                     ; //=8'h73
   reg signed [  3:  0] W0245                     ; //=4'hf
   reg signed [  2:  0] W0246                     ; //=3'h7
   reg signed [ 74:  0] W0247 /*verilator public*/; //=75'h0000000000000000000
   reg signed [ 27:  0] W0248                     ; //=28'h0000000
   reg        [ 42:  0] W0249 /*verilator public*/; //=43'h7ffffffffff
   reg signed [ 92:  0] W0250                     ; //=93'h000000000000000000000000
   reg        [ 54:  0] W0251                     ; //=55'h00000000000000
   reg        [ 95:  0] W0252                     ; //=96'h000000000000000000000000
   reg signed [ 38:  0] W0253                     ; //=39'h005f38482c
   reg signed [ 78:  0] W0254                     ; //=79'h7fff87182181ffffffff
   reg        [126:  0] W0255 /*verilator public*/; //=127'h00000000000000000000000000000000
   reg signed [ 77:  0] W0256                     ; //=78'h000200000002951e42d6
   reg        [  0:  0] W0257                     ; //=1'h1
   reg        [112:  0] W0258                     ; //=113'h00000000000000000000000000000
   reg signed [ 80:  0] W0259 /*verilator public*/; //=81'h1ffffffffffffffffffff
   reg        [ 35:  0] W0260                     ; //=36'h000000000
   reg        [102:  0] W0261 /*verilator public*/; //=103'h00000000000000000000000000
   reg signed [113:  0] W0262                     ; //=114'h00000000000000000000000000000
   reg        [ 47:  0] W0263                     ; //=48'h000000000000
   reg signed [127:  0] W0264 /*verilator public*/; //=128'h00000000000000000000000000000000
   reg signed [ 34:  0] W0265                     ; //=35'h000000000
   reg signed [ 30:  0] W0266 /*verilator public*/; //=31'h7fffffff
   reg        [ 90:  0] W0267                     ; //=91'h73a41afffffffffffffffff
   reg signed [ 50:  0] W0268                     ; //=51'h00000e748356c
   reg signed [127:  0] W0269                     ; //=128'hffffffffffffffffffffffffffffffff
   reg signed [ 18:  0] W0270                     ; //=19'h00000
   reg signed [ 53:  0] W0271                     ; //=54'h00000000000001
   reg        [ 82:  0] W0272 /*verilator public*/; //=83'h51274ffffffffffffffff
   reg        [ 34:  0] W0273                     ; //=35'h000000001
   reg        [ 16:  0] W0274 /*verilator public*/; //=17'h00000
   reg signed [ 66:  0] W0275 /*verilator public*/; //=67'h00000000000000000
   reg signed [102:  0] W0276 /*verilator public*/; //=103'h00000000000000000000000001
   reg        [  5:  0] W0277                     ; //=6'h3f
   reg signed [  9:  0] W0278                     ; //=10'h3ff
   reg signed [122:  0] W0279 /*verilator public*/; //=123'h0000000feefe6b4ffffffffc7107e4a
   reg        [  0:  0] W0280 /*verilator public*/; //=1'h0
   reg        [ 49:  0] W0281                     ; //=50'h0000000000000
   reg        [ 49:  0] W0282 /*verilator public*/; //=50'h0000000000000
   reg        [ 78:  0] W0283                     ; //=79'h7fffffffffffffffff84
   reg        [127:  0] W0284                     ; //=128'hfffffffffffffffffffffffe101dee12
   reg        [ 94:  0] W0285                     ; //=95'h7fffffffffffffffffffffff
   reg signed [ 66:  0] W0286 /*verilator public*/; //=67'h00000000000000000
   reg        [  0:  0] W0287                     ; //=1'h0
   reg signed [  1:  0] W0288                     ; //=2'h3
   reg signed [124:  0] W0289                     ; //=125'h00000000000000000000000000000000
   reg        [112:  0] W0290 /*verilator public*/; //=113'h00000000000000006d1262eca71c0
   reg signed [120:  0] W0291                     ; //=121'h1906da100000001ffffffff00000000
   reg signed [120:  0] W0292 /*verilator public*/; //=121'h1906da100000001ffffffff00000000
   reg        [120:  0] W0293 /*verilator public*/; //=121'h0000000000000001fffffffffc05c47
   reg signed [127:  0] W0294                     ; //=128'h0000000000000000fffffffffe02e239
   reg signed [127:  0] W0295 /*verilator public*/; //=128'h0000000100000000d0ed7551a8e8b0f8
   reg        [121:  0] W0296                     ; //=122'h3ffffffffffffffffffffffffffffff
   reg        [ 58:  0] W0297                     ; //=59'h7ffffffffffffff
   reg signed [ 78:  0] W0298                     ; //=79'h7fffffffffffffffffff
   reg signed [110:  0] W0299 /*verilator public*/; //=111'h7fffffffffffffffffffffffffff
   reg signed [ 54:  0] W0300                     ; //=55'h00000000000000
   reg signed [ 26:  0] W0301                     ; //=27'h7ffffff
   reg signed [ 17:  0] W0302                     ; //=18'h00002
   reg signed [  6:  0] W0303                     ; //=7'h7f
   reg        [110:  0] W0304                     ; //=111'h0000000000000000000000000000
   reg        [ 96:  0] W0305                     ; //=97'h0000000000000000000374acf
   reg signed [115:  0] W0306 /*verilator public*/; //=116'h000004a144132ffffffffffffffff
   reg        [ 19:  0] W0307                     ; //=20'h00000
   reg signed [ 22:  0] W0308 /*verilator public*/; //=23'h283d11
   reg        [ 85:  0] W0309                     ; //=86'h0000000000000000000000
   reg signed [127:  0] W0310                     ; //=128'hffffffffffffffffffffffffffffffff
   reg signed [127:  0] W0311                     ; //=128'hffffffffffffffffffffffffffffffff
   reg        [ 53:  0] W0312 /*verilator public*/; //=54'h00000000000000
   reg signed [110:  0] W0313                     ; //=111'h0000000000000000000000000000
   reg signed [110:  0] W0314                     ; //=111'h0000000000000000000000000000
   reg signed [110:  0] W0315                     ; //=111'h0000000000000000000000000000
   reg signed [127:  0] W0316 /*verilator public*/; //=128'hffffffffffffffffffffffffffffffff
   reg signed [ 80:  0] W0317                     ; //=81'h13544d664fd48350489be
   reg signed [ 80:  0] W0318                     ; //=81'h000006ff7e650350489be
	//============================================================
   always @(check) begin : Block1
	W0003 = 128'shffffffffffffffffffffffffffffffff;
	W0002 = (4'hf << {1'h1,2'h3});
	W0001 = W0003;
	if (96'sh0 != 96'sh0) if (check) $stop;
	if (W0001[W0002+:96] != 96'hffffffffffffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block2
	if ((~ {4'h0,((59'h0 >> 7'h7f) ^ (1'h0 ? 59'h0 : 59'h7ffffffffffffff))}) != 63'h7800000000000000) if (check) $stop;
	if ((((((100'shfffffffff17d4750300000000 >>> 8'sh0) & (100'sh000000000ffffffff68138f72 >>> 8'shff)))==100'h0 ? 100'sh0:(100'sh14bb5d8e3ffffffffeda1130c / ((100'shfffffffff17d4750300000000 >>> 8'sh0) & (100'sh000000000ffffffff68138f72 >>> 8'shff)))) >>> (- ((8'shb3 >>> 4'sh1) <<< 4'sh0))) != 100'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0007 <= 95'sh1feb10faffffffff00000000;
   end
   always @(posedge clk) begin
	W0006 <= 36'sh000000001;
   end
   always @(posedge clk) begin
	W0005 <= ((3'h7)==3'h0 ? 3'h0:(3'h1 % 3'h7));
   end
   always @(posedge clk) begin
	W0004 <= 119'h2f54d600000000ffffffff00000000;
   end
   always @(posedge clk) begin
	if (W0004[5'h0+:64] != 64'hffffffff00000000) if (check) $stop;
	if ($unsigned((W0005[2+:1] ? W0006[35:34] : {1'h0,W0007[6'h3f]})) != 2'h1) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block4
	W0008 = 61'h1fffffffffffffff;
	if (2'sh3 != 2'sh3) if (check) $stop;
	if ((~ ((W0008[60:60])==1'h0 ? 1'h0:((((65'sh0ffffffffffffffff)==65'h0 ? 65'sh0:(65'sh0 % 65'sh0ffffffffffffffff)) !== (65'sh00000000000000001 >>> 8'shff)) / W0008[60:60]))) != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0013 <= 109'h1fffffffffffffffffffffffffff;
   end
   always @(posedge clk) begin
	W0012 <= W0013;
   end
   always @(posedge clk) begin
	W0011 <= W0012[108:102];
   end
   always @(posedge clk) begin
	W0010 <= ((63'sh7fffffffffffffff)==63'h0 ? 63'sh0:(63'sh7fffffffffffffff / 63'sh7fffffffffffffff));
   end
   always @(posedge clk) begin
	W0009 <= ((102'sh3f3ec596b700000000d12d2796)==102'h0 ? 102'sh0:(102'sh0 % 102'sh3f3ec596b700000000d12d2796));
   end
   always @(posedge clk) begin
	if ((((~ W0009))==102'h0 ? 102'sh0:(102'sh00ffffffffffffffff38390476 % (~ W0009))) != 102'sh0) if (check) $stop;
	if ((((61'h0000000180c90692)==61'h0 ? 61'h0:(W0010[2+:61] / 61'h0000000180c90692)) >> W0011) != 61'h0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block6
	W0017 = (($unsigned(1'h1) ? (32'shffffffff >>> 6'sh0) : (32'shffffffff | 32'shffffffff)) + ((32'shca1cfecf <<< 6'sh3f) <<< 6'sh0a));
	W0016 = 88'sh0;
	W0015 = 8'sh0;
	W0014 = (((~ W0016[87:21]))==67'h0 ? 67'h0:({W0015,59'sh0} % (~ W0016[87:21])));
	if (W0014[62-:63] != 63'h0) if (check) $stop;
	if (W0017 != 32'shffffffff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0020 <= 97'sh1ffffffffffffffffffffffff;
   end
   always @(posedge clk) begin
	W0019 <= (97'sh000000001abf37a3000000000 + 97'sh0000000000000000000000001);
   end
   always @(posedge clk) begin
	W0018 <= ((((124'shfffffffffffffffffffffffffffffff)==124'h0 ? 124'sh0:(124'shfffffffffffffffffffffffffffffff / 124'shfffffffffffffffffffffffffffffff)) >>> 8'shff) >>> 8'sh68);
   end
   always @(posedge clk) begin
	if (W0018[123:123] != 1'h0) if (check) $stop;
	if (((W0020)==97'h0 ? 97'sh0:(((W0019)==97'h0 ? 97'sh0:((~ 97'sh0ffffffffffffffff648b6e1f) % W0019)) / W0020)) != 97'sh00000000119d226becb67d8c4) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0022 <= 123'sh7ffffffbce03e2bdb14609fe7e28b41;
   end
   always @(posedge clk) begin
	W0021 <= 126'sh3fffffffffffffffffffffffffffffff;
   end
   always @(posedge clk) begin
	if (W0021[125:125] != 1'h1) if (check) $stop;
	if (W0022[94-:95] != 95'h3ce03e2bdb14609fe7e28b41) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block9
	if (102'sh3fffffffffffffffffffffffff != 102'sh3fffffffffffffffffffffffff) if (check) $stop;
	if (9'h1ff != 9'h1ff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0030 <= 95'sh3691dbd700000000ffffffff;
   end
   always @(posedge clk) begin
	W0029 <= (((95'sh7fffffffffffffffffffffff <<< 8'shff))==95'h0 ? 95'sh0:(W0030 / (95'sh7fffffffffffffffffffffff <<< 8'shff)));
   end
   always @(posedge clk) begin
	W0028 <= (- 39'sh7fa0c7b7d4);
   end
   always @(posedge clk) begin
	W0027 <= (7'sh7f >>> 4'sh1);
   end
   always @(posedge clk) begin
	W0026 <= W0028;
   end
   always @(posedge clk) begin
	W0025 <= W0029[94:20];
   end
   always @(posedge clk) begin
	W0024 <= ((~ 84'shf099500000001cf74c284) - 84'shfffffffffffffffffffff);
   end
   always @(posedge clk) begin
	W0023 <= (~ 84'shfffffffffffff1e016f6b);
   end
   always @(posedge clk) begin
	if (((W0024)==84'h0 ? 84'sh0:($signed(W0023) % W0024)) != 84'sh0000000000000e1fe9094) if (check) $stop;
	if (W0025[W0026[W0027[2+:5]+:6]+:2] != 2'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0032 <= (64'sh00000001ffffffff * 64'shffffffffffffffff);
   end
   always @(posedge clk) begin
	W0031 <= (W0032 >>> ((1'h0 ? 7'sh4d : 7'sh27) & (~ 7'sh7f)));
   end
   always @(posedge clk) begin
	if (W0031 != 64'shfffffffe00000001) if (check) $stop;
	if (2'sh1 != 2'sh1) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block12
	W0033 = 32'hffffffff;
	if (((((~ $signed(2'h0)) >>> (2'sh0 >>> (2'sh1 >>> 2'sh3))))==2'h0 ? 2'sh0:(2'sh3 % ((~ $signed(2'h0)) >>> (2'sh0 >>> (2'sh1 >>> 2'sh3))))) != 2'sh0) if (check) $stop;
	if (((W0033[31:31])==1'h0 ? 1'h0:(1'h1 % W0033[31:31])) != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(check or W0009 or W0017) begin : Block13
   end
   always @(posedge clk) begin : Block13Check
	if (W0009 != 102'sh0) if (check) $stop;
	if (W0017 != 32'shffffffff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0038 <= ((3'sh0)==3'h0 ? 3'sh0:(3'sh7 % 3'sh0));
   end
   always @(posedge clk) begin
	W0037 <= 31'sh7fffffff;
   end
   always @(posedge clk) begin
	W0036 <= (95'h7fffffffffffffffffffffff - 95'h0000000023324557404ae610);
   end
   always @(posedge clk) begin
	W0035 <= (90'sh3ffffff5165d0f4ffffffff ^ 90'sh3ffffffffffffffffffffff);
   end
   always @(posedge clk) begin
	W0034 <= W0036;
   end
   always @(posedge clk) begin
	if (((60'sh000000000000001 === (((1'h0 ? 60'sh0 : 60'sh0))==60'h0 ? 60'sh0:(((60'sh000000000000001)==60'h0 ? 60'sh0:(60'shff9e16800000000 % 60'sh000000000000001)) / (1'h0 ? 60'sh0 : 60'sh0)))) ? W0034[W0035[89:84]+:1] : (~ (W0037 && W0032))) != 1'h0) if (check) $stop;
	if (W0038[2:2] != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if ((1'h1 ? 72'shff55c5414cc8a8bf33 : 72'shffffffffffffffffff) != 72'shff55c5414cc8a8bf33) if (check) $stop;
	if ((110'sh0000000000000000000000000001 >>> ((8'shff)==8'h0 ? 8'sh0:(($signed(8'sh0) >>> (4'shf <<< 3'sh7)) % 8'shff))) != 110'sh0000000000000000000000000001) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0040 <= ((4'sh0)==4'h0 ? 4'sh0:(4'sh1 % 4'sh0));
   end
   always @(posedge clk) begin
	W0039 <= (67'sh200000001fc7de7a7 <<< ((W0015)==8'h0 ? 8'sh0:(W0015 / W0015)));
   end
   always @(posedge clk) begin
	if (W0039[3+:64] != 64'h400000003f8fbcf4) if (check) $stop;
	if ((((W0030)==95'h0 ? 95'sh0:(W0030 % W0030)) <<< (W0015 >>> W0040)) != 95'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (1'h0 != 1'h0) if (check) $stop;
	if ((28'sh0000001 <<< ((((6'sh0 >>> 4'shf))==6'h0 ? 6'sh0:((6'sh0 >>> 4'sh1) / (6'sh0 >>> 4'shf))) | (6'sh3f <<< ((4'sh0)==4'h0 ? 4'sh0:(4'shf / 4'sh0))))) != 28'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (W0037 != 31'sh7fffffff) if (check) $stop;
	if (60'h0 != 60'h0) if (check) $stop;
   end
	//============================================================
   always @(check or W0037) begin : Block19
	W0043 = 99'sh7ffffffffffffffffffffffff;
	W0042 = 7'sh7f;
	W0041 = (31'sh7fffffff - W0037);
	if ((~ W0041) != 31'sh7fffffff) if (check) $stop;
	if ((((((44'sh0 >>> 7'sh01) >>> W0042) >>> (W0043[27-:1] ? ((7'sh01)==7'h0 ? 7'sh0:(7'sh0 % 7'sh01)) : (7'sh0 >>> 4'shf))))==44'h0 ? 44'sh0:((((1'h1 ? 44'sh0 : 44'sh928eff62598) >>> 7'sh7f) <<< (7'sh01 >>> (4'shf >>> 3'sh0))) % (((44'sh0 >>> 7'sh01) >>> W0042) >>> (W0043[27-:1] ? ((7'sh01)==7'h0 ? 7'sh0:(7'sh0 % 7'sh01)) : (7'sh0 >>> 4'shf))))) != 44'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0046 <= (85'h1fffffffffffffffffffff << 8'hd9);
   end
   always @(posedge clk) begin
	W0045 <= (107'h0 << 8'hff);
   end
   always @(posedge clk) begin
	W0044 <= ((W0046)==85'h0 ? 85'h0:(W0045[106:22] % W0046));
   end
   always @(posedge clk) begin
	if (($signed((((5'h1f << 4'hf))==5'h0 ? 5'h0:(((5'h1f)==5'h0 ? 5'h0:(5'h0 / 5'h1f)) % (5'h1f << 4'hf)))) <<< (W0040 >>> (((3'sh7)==3'h0 ? 3'sh0:(3'sh0 % 3'sh7)) >>> (3'sh7 >>> 3'sh0)))) != 5'sh0) if (check) $stop;
	if (W0044[84:83] != 2'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (42'h0 != 42'h0) if (check) $stop;
	if (1'h1 != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0047 <= (96'shffffffffffffffffffffffff <<< W0015);
   end
   always @(posedge clk) begin
	if (W0047 != 96'shffffffffffffffffffffffff) if (check) $stop;
	if (1'h0 != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0049 <= ((((51'sh7ffffffffffff)==51'h0 ? 51'sh0:((51'sh7ffffffffffff >>> 7'sh54) % 51'sh7ffffffffffff)))==51'h0 ? 51'sh0:(51'sh7ffffffffffff % ((51'sh7ffffffffffff)==51'h0 ? 51'sh0:((51'sh7ffffffffffff >>> 7'sh54) % 51'sh7ffffffffffff))));
   end
   always @(posedge clk) begin
	W0048 <= 63'h00000001bf003b47;
   end
   always @(posedge clk) begin
	if (W0048[62:53] != 10'h0) if (check) $stop;
	if (W0049[50:50] != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0051 <= (108'sh0170f5f330fffffffff5d6adc0c + 108'shfffffffffffffffffffffffffff);
   end
   always @(posedge clk) begin
	W0050 <= (((1'h0 ? 108'sh0 : 108'sh0) <<< ((8'sh0)==8'h0 ? 8'sh0:(8'sh0 % 8'sh0))) | W0051);
   end
   always @(posedge clk) begin
	if (W0050[107:40] != 68'h0170f5f330fffffff) if (check) $stop;
	if (31'h7fffffff != 31'h7fffffff) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block25
	W0054 = (2'sh3 - 2'sh3);
	W0053 = (2'sh0 >>> 2'sh0);
	W0052 = (((2'sh0)==2'h0 ? 2'sh0:(2'sh3 / 2'sh0)) ^ (2'sh3 <<< 2'sh2));
	if ((((W0053 >>> (((2'sh3)==2'h0 ? 2'sh0:(2'sh0 / 2'sh3)) <<< ((2'sh3)==2'h0 ? 2'sh0:(2'sh0 / 2'sh3)))))==2'h0 ? 2'sh0:(W0052 / (W0053 >>> (((2'sh3)==2'h0 ? 2'sh0:(2'sh0 / 2'sh3)) <<< ((2'sh3)==2'h0 ? 2'sh0:(2'sh0 / 2'sh3)))))) != 2'sh0) if (check) $stop;
	if (((2'sh3)==2'h0 ? 2'sh0:((W0054 <<< (2'sh0 <<< (2'sh1 >>> 2'sh0))) / 2'sh3)) != 2'sh0) if (check) $stop;
   end
	//============================================================
   always @(check or W0052) begin : Block26
	if (99'sh153fb34be2a39f49d00000000 != 99'sh153fb34be2a39f49d00000000) if (check) $stop;
	if ((W0052 | 2'sh0) != 2'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0057 <= (- 53'h156230ffffffff);
   end
   always @(posedge clk) begin
	W0056 <= 20'sh0;
   end
   always @(posedge clk) begin
	W0055 <= 71'sh0;
   end
   always @(posedge clk) begin
	if ((W0055[W0056[19:14]+:1] | (& W0057[52:52])) != 1'h0) if (check) $stop;
	if (((((40'sh0 <<< 7'sh7f) <<< ((((7'sh51)==7'h0 ? 7'sh0:(7'sh7f % 7'sh51)))==7'h0 ? 7'sh0:(((7'sh7f)==7'h0 ? 7'sh0:(7'sh7f % 7'sh7f)) / ((7'sh51)==7'h0 ? 7'sh0:(7'sh7f % 7'sh51))))))==40'h0 ? 40'sh0:(40'shffffffffff / ((40'sh0 <<< 7'sh7f) <<< ((((7'sh51)==7'h0 ? 7'sh0:(7'sh7f % 7'sh51)))==7'h0 ? 7'sh0:(((7'sh7f)==7'h0 ? 7'sh0:(7'sh7f % 7'sh7f)) / ((7'sh51)==7'h0 ? 7'sh0:(7'sh7f % 7'sh51))))))) != 40'sh0) if (check) $stop;
   end
	//============================================================
   always @(check or W0032) begin : Block28
	W0060 = 128'h0;
	W0059 = $signed(85'sh1fffffffffffffc422fb6e);
	W0058 = ((W0060[4'h5+:99])==99'h0 ? 99'h0:(99'h7ffffffffffffffffffffffff % W0060[4'h5+:99]));
   end
   always @(posedge clk) begin : Block28Check
	if ((~ W0058[W0059[84:80]+:64]) != 64'hffffffffffffffff) if (check) $stop;
	if (W0032 != 64'shfffffffe00000001) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0064 <= 25'sh1ffffff;
   end
   always @(posedge clk) begin
	W0063 <= 28'sh0;
   end
   always @(posedge clk) begin
	W0062 <= 61'sh1fffffffffffffff;
   end
   always @(posedge clk) begin
	W0061 <= W0062[60:60];
   end
   always @(posedge clk) begin
	if (W0061 != 1'h1) if (check) $stop;
	if ((W0063[27:27] & W0064[24:24]) != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(check or W0042) begin : Block30
	W0068 = (15'sh0 + 15'sh0);
	W0067 = 51'h0;
	W0066 = (8'sh1e >>> 4'shf);
	W0065 = (128'shffffffffffffffffffffffffffffffff <<< 8'sh0);
   end
   always @(posedge clk) begin : Block30Check
	if ((({(45'sh1fffffffffff >>> W0042),W0067})==96'h0 ? 96'h0:(W0065[W0066[7:4]+:96] / {(45'sh1fffffffffff >>> W0042),W0067})) != 96'h000000000000000000000001) if (check) $stop;
	if (((((~ (15'sh0001 >>> 5'sh1f)))==15'h0 ? 15'sh0:(W0068 % (~ (15'sh0001 >>> 5'sh1f)))) >>> 5'sh1f) != 15'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0072 <= ((126'sh3fffffffffffffffffffffffffffffff)==126'h0 ? 126'sh0:(126'sh00000000000000000000000000000001 % 126'sh3fffffffffffffffffffffffffffffff));
   end
   always @(posedge clk) begin
	W0071 <= 123'h0;
   end
   always @(posedge clk) begin
	W0070 <= W0071;
   end
   always @(posedge clk) begin
	W0069 <= (W0070 + W0072[125:3]);
   end
   always @(posedge clk) begin
	if (21'h0 != 21'h0) if (check) $stop;
	if (W0069 != 123'h0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block32
	W0077 = 99'sh7ffffffffffffffffffffffff;
	W0076 = (126'h3fffffff000000015e4ef77c00000000 >> W0077[61-:8]);
	W0075 = W0076[125:0];
	W0074 = ((((39'sh7fffffffff)==39'h0 ? 39'sh0:(39'sh0 / 39'sh7fffffffff)))==39'h0 ? 39'sh0:(((39'sh0)==39'h0 ? 39'sh0:(39'sh7f2a25b834 % 39'sh0)) / ((39'sh7fffffffff)==39'h0 ? 39'sh0:(39'sh0 / 39'sh7fffffffff))));
	W0073 = 51'sh7ffffffffffff;
   end
   always @(posedge clk) begin : Block32Check
	if (W0073[W0074[31-:5]+:1] != 1'h1) if (check) $stop;
	if (W0075[125:30] != 96'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0078 <= {4{((1'h0 ? 6'sh06 : 6'sh01) | (6'sh3f >>> 4'shb))}};
   end
   always @(posedge clk) begin
	if (W0078[23:23] != 1'h1) if (check) $stop;
	if (((16'shffff <= ((16'sh0042 >>> 5'sh0) >>> ((5'sh0)==5'h0 ? 5'sh0:(5'sh1f / 5'sh0)))) >> ((^~ (41'h0 | 41'h1ff2efa1bb2)) === ({7'h0,111'h767cffffffff3d032af100000000} || (~ 10'sh0)))) != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0081 <= 111'sh5d8cffffffff9b20638fffffffff;
   end
   always @(posedge clk) begin
	W0080 <= 8'h0;
   end
   always @(posedge clk) begin
	W0079 <= ((({64'sh1e9f5381b93a757b,62'sh0} << W0080))==126'h0 ? 126'h0:($unsigned((126'sh00000000000000000000000000000001 & 126'sh0)) % ({64'sh1e9f5381b93a757b,62'sh0} << W0080)));
   end
   always @(posedge clk) begin
	if (W0079 != 126'h0) if (check) $stop;
	if (W0081[110:79] != 32'hbb19ffff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0082 <= 14'sh0;
   end
   always @(posedge clk) begin
	if ((! W0082) != 1'h1) if (check) $stop;
	if (113'h00000ffffffff07a5ea017b37c2ff != 113'h00000ffffffff07a5ea017b37c2ff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0084 <= 6'sh30;
   end
   always @(posedge clk) begin
	W0083 <= 32'sh0;
   end
   always @(posedge clk) begin
	if (((W0047)==96'h0 ? 96'sh0:(W0047 % W0047)) != 96'sh0) if (check) $stop;
	if ((((((W0017 >>> W0084))==32'h0 ? 32'sh0:(W0083 % (W0017 >>> W0084))))==32'h0 ? 32'sh0:((W0017 | ((((32'sh0)==32'h0 ? 32'sh0:(32'sh0 % 32'sh0)))==32'h0 ? 32'sh0:((~ 32'sha60d289a) / ((32'sh0)==32'h0 ? 32'sh0:(32'sh0 % 32'sh0))))) / (((W0017 >>> W0084))==32'h0 ? 32'sh0:(W0083 % (W0017 >>> W0084))))) != 32'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if ((((((17'sh1ffff)==17'h0 ? 17'sh0:((~ 17'sh0) % 17'sh1ffff)) <<< 6'sh3f))==17'h0 ? 17'sh0:(17'sh0973d / (((17'sh1ffff)==17'h0 ? 17'sh0:((~ 17'sh0) % 17'sh1ffff)) <<< 6'sh3f))) != 17'sh0) if (check) $stop;
	if (15'sh7fff != 15'sh7fff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0090 <= (((6'sh3f)==6'h0 ? 6'sh0:(6'sh0 / 6'sh3f)) + 6'sh1b);
   end
   always @(posedge clk) begin
	W0089 <= 79'sh0;
   end
   always @(posedge clk) begin
	W0088 <= W0089[78:11];
   end
   always @(posedge clk) begin
	W0087 <= 26'sh0000001;
   end
   always @(posedge clk) begin
	W0086 <= (51'sh0 & 51'sh0);
   end
   always @(posedge clk) begin
	W0085 <= ((90'sh3ffffffffffffffffffffff <<< 8'sh0) >>> (1'h1 ? 8'shff : 8'sh0));
   end
   always @(posedge clk) begin
	if (((((W0088[67:66])==2'h0 ? 2'h0:(W0086[W0087[25:21]+:2] % W0088[67:66])))==2'h0 ? 2'h0:(W0085[89:88] / ((W0088[67:66])==2'h0 ? 2'h0:(W0086[W0087[25:21]+:2] % W0088[67:66])))) != 2'h0) if (check) $stop;
	if ((18'sh3ffff >>> W0090) != 18'sh3ffff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (72'shffffffffffffffffff != 72'shffffffffffffffffff) if (check) $stop;
	if (98'sh000000001cf98bdd8ed1bf345 != 98'sh000000001cf98bdd8ed1bf345) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0092 <= 78'sh3fffffffffffffffffff;
   end
   always @(posedge clk) begin
	W0091 <= (W0092 >>> (8'sh0 <<< 4'sh0));
   end
   always @(posedge clk) begin
	if (((W0091)==78'h0 ? 78'sh0:((((((78'sh0)==78'h0 ? 78'sh0:(78'sh3fffffffffff64616519 / 78'sh0)) >>> W0015))==78'h0 ? 78'sh0:((78'sh3fffffffffffffffffff <<< ((8'sh01)==8'h0 ? 8'sh0:(8'shff % 8'sh01))) / (((78'sh0)==78'h0 ? 78'sh0:(78'sh3fffffffffff64616519 / 78'sh0)) >>> W0015))) / W0091)) != 78'sh0) if (check) $stop;
	if ((- ($signed(((49'sh0)==49'h0 ? 49'sh0:(49'sh1ffffffffffff % 49'sh0))) >>> 7'sh6b)) != 49'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0093 <= W0003;
   end
   always @(posedge clk) begin
	if (W0093[99-:95] != 95'h7fffffffffffffffffffffff) if (check) $stop;
	if (W0047 != 96'shffffffffffffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block42
	W0095 = 19'sh7ffff;
	W0094 = (((127'sh0 >>> 8'sh0))==127'h0 ? 127'sh0:(((127'sh7fffffffffffffffffffffffffffffff)==127'h0 ? 127'sh0:(127'sh00000000000000000000000000000001 / 127'sh7fffffffffffffffffffffffffffffff)) % (127'sh0 >>> 8'sh0)));
	if (106'sh3ffc3b5c523ffffffffffffffff != 106'sh3ffc3b5c523ffffffffffffffff) if (check) $stop;
	if ((W0094[126:15] << W0095[12-:8]) != 112'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0098 <= W0003;
   end
   always @(posedge clk) begin
	W0097 <= W0003;
   end
   always @(posedge clk) begin
	W0096 <= W0015;
   end
   always @(posedge clk) begin
	if ((((80'shffff41044a6b00000001 >>> (8'shff >>> 4'sh0)) | (~ 80'sh0)) >>> W0096) != 80'shffffffffffffffffffff) if (check) $stop;
	if (((W0098[4'h0+:97])==97'h0 ? 97'h0:(((W0097[4'h1+:97])==97'h0 ? 97'h0:({1{(97'sh0 <<< 8'shff)}} % W0097[4'h1+:97])) / W0098[4'h0+:97])) != 97'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0100 <= (1'h1 ? 20'shfffff : 20'sh0);
   end
   always @(posedge clk) begin
	W0099 <= (((20'sh0 >>> (6'sh3f >>> 4'sh0)))==20'h0 ? 20'sh0:(W0100 / (20'sh0 >>> (6'sh3f >>> 4'sh0))));
   end
   always @(posedge clk) begin
	if ((- 86'sh0) != 86'sh0) if (check) $stop;
	if (W0099 != 20'sh0) if (check) $stop;
   end
	//============================================================
   always @(check or W0061) begin : Block45
	W0101 = ((75'sh7ff7e019ac646679f3d >>> 8'sh0) ^ 75'sh0);
   end
   always @(posedge clk) begin : Block45Check
	if ($signed(W0101[74:16]) != 59'sh7ff7e019ac64667) if (check) $stop;
	if (W0061 != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(check or W0096) begin : Block46
	W0104 = (122'sh3ffffff000000010000000000000001 >>> 8'shff);
	W0103 = (W0104 >>> W0096);
	W0102 = ((((86'sh0 >>> 8'sh01) | 86'sh16da685016495100000000))==86'h0 ? 86'sh0:(((86'sh3fffffffffffffffffffff >>> 8'sh01) <<< (8'sh0 >>> 4'sh1)) % ((86'sh0 >>> 8'sh01) | 86'sh16da685016495100000000)));
	if (W0102 != 86'sh3fffffffffffffffffffff) if (check) $stop;
	if (W0103[121:91] != 31'h7fffffff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if ((53'sh000000391b7da7 ^ (~ ((53'sh1fffffffffffff)==53'h0 ? 53'sh0:((1'h0 ? 53'sh000000ffffffff : 53'sh1fffffffffffff) % 53'sh1fffffffffffff)))) != 53'sh1fffffc6e48258) if (check) $stop;
	if ((~ 5'h0) != 5'h1f) if (check) $stop;
   end
	//============================================================
   always @(check or W0031 or W0096) begin : Block48
	W0107 = 89'sh1ffffff04b841e1ffffffff;
	W0106 = ((89'sh0 >>> W0096) - W0107);
	W0105 = (4'shf & 4'sh0);
	if (((W0031 >>> (((7'sh7f)==7'h0 ? 7'sh0:(7'sh0 / 7'sh7f)) >>> 4'shf)) >>> (((7'sh0 & 7'sh7f) | (7'sh0 <<< 4'sh4)) <<< W0105)) != 64'shfffffffe00000001) if (check) $stop;
	if (W0106 != 89'sh0000000fb47be1e00000001) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (((48'sh00009b021b77)==48'h0 ? 48'sh0:(((48'shc4c800000001)==48'h0 ? 48'sh0:(48'sh30853054aa34 / 48'shc4c800000001)) / 48'sh00009b021b77)) != 48'sh0) if (check) $stop;
	if ((71'sh0 ^ 71'sh0) != 71'sh0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block50
	W0109 = (((67'sh7ffffffffffffffff)==67'h0 ? 67'sh0:(67'sh7ffffffffffffffff / 67'sh7ffffffffffffffff)) * (67'sh0ffffffff29ed52ab >>> 8'shff));
	W0108 = W0109;
	if (W0108[1'h0+:63] != 63'h0) if (check) $stop;
	if (29'sh0 != 29'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0110 <= $signed(61'h0);
   end
   always @(posedge clk) begin
	if (W0110 != 61'sh0) if (check) $stop;
	if (((115'sh7ffffffffffffffffffff00000000 >>> (((8'sh01)==8'h0 ? 8'sh0:(8'shff % 8'sh01)) <<< W0040)) >>> 8'shff) != 115'sh7ffffffffffffffffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(check or W0061) begin : Block52
	W0113 = 40'h0;
	W0112 = $unsigned(W0113);
	W0111 = 7'sh01;
   end
   always @(posedge clk) begin : Block52Check
	if ((((~ ((63'sh000000001976eaa4 >>> 7'sh7c) >>> 7'sh01)))==63'h0 ? 63'sh0:((63'sh0 & ((1'h1 ? 63'sh0 : 63'sh0) >>> W0111)) % (~ ((63'sh000000001976eaa4 >>> 7'sh7c) >>> 7'sh01)))) != 63'sh0) if (check) $stop;
	if ((W0061 >> W0112[39:39]) != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(check or W0080 or W0083) begin : Block53
	W0118 = 88'sh0;
	W0117 = W0118;
	W0116 = (81'h000000000000000000001 << 8'h0);
	W0115 = 79'sh0001ffffffff00000000;
	W0114 = W0115;
	if (W0083 != 32'sh0) if (check) $stop;
	if ((((W0117[87:13] << W0080))==75'h0 ? 75'h0:(((W0116[80:6])==75'h0 ? 75'h0:(W0114[78:4] / W0116[80:6])) / (W0117[87:13] << W0080))) != 75'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0122 <= (38'sh3fffffffff + 38'sh0000000001);
   end
   always @(posedge clk) begin
	W0121 <= 40'h0;
   end
   always @(posedge clk) begin
	W0120 <= W0121[39:39];
   end
   always @(posedge clk) begin
	W0119 <= (99'h1ffffffffb8784d1000000001 >> 8'h01);
   end
   always @(posedge clk) begin
	if (((W0119[27-:1] <  W0120) ? ((~ (63'sh7fffffffffffffff <<< 7'sh0)) >>> W0111) : (~ (63'sh0 >>> (7'sh7f >>> 4'shf)))) != 63'sh7fffffffffffffff) if (check) $stop;
	if (((~ W0122) <<< 7'sh65) != 38'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0123 <= 46'sh0;
   end
   always @(posedge clk) begin
	if ((((((1'h0 ? 46'sh0 : 46'sh353300000000) >>> (1'h0 ? 7'sh0 : 7'sh0)) >>> $signed(W0111)))==46'h0 ? 46'sh0:((((W0123 >>> W0042))==46'h0 ? 46'sh0:(($signed(46'sh0) >>> W0111) % (W0123 >>> W0042))) % (((1'h0 ? 46'sh0 : 46'sh353300000000) >>> (1'h0 ? 7'sh0 : 7'sh0)) >>> $signed(W0111)))) != 46'sh0) if (check) $stop;
	if (((1'h1)==1'h0 ? 1'h0:(1'h0 % 1'h1)) != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0125 <= W0080;
   end
   always @(posedge clk) begin
	W0124 <= {1{71'sh7fffffffffffffffff}};
   end
   always @(posedge clk) begin
	if (84'sh00000ffffffff00000000 != 84'sh00000ffffffff00000000) if (check) $stop;
	if ((((W0124 >> W0125))==71'h0 ? 71'h0:(((71'h000000000000000001)==71'h0 ? 71'h0:(71'h05ffffffff00000000 % 71'h000000000000000001)) % (W0124 >> W0125))) != 71'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0127 <= (76'sh0 - 76'sh0000000000000000001);
   end
   always @(posedge clk) begin
	W0126 <= (83'sh7ffff00000000397f927d >>> 8'sh0);
   end
   always @(posedge clk) begin
	if ((1'h1 ? (^ W0126[82:20]) : 1'h0) != 1'h0) if (check) $stop;
	if (((W0127 ^ (((76'sh0000000000000000001 >>> 8'sh69))==76'h0 ? 76'sh0:(76'shd6f3f197a9e00000000 / (76'sh0000000000000000001 >>> 8'sh69)))) >>> (8'shff | W0096)) != 76'shfffffffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0130 <= 128'shffffffffffffffffffffffffffffffff;
   end
   always @(posedge clk) begin
	W0129 <= 52'hfffffffffffff;
   end
   always @(posedge clk) begin
	W0128 <= W0068;
   end
   always @(posedge clk) begin
	if (W0128[12-:13] != 13'h0) if (check) $stop;
	if ({((38'h1d69b1ac3b)==38'h0 ? 38'h0:(((W0130[6'h0+:38])==38'h0 ? 38'h0:(W0129[51:14] / W0130[6'h0+:38])) % 38'h1d69b1ac3b)),26'h0} != 64'h0000000004000000) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0132 <= (~ 126'sh01165f8a0000000010f0cce7a72797f4);
   end
   always @(posedge clk) begin
	W0131 <= 67'sh00000000000000001;
   end
   always @(posedge clk) begin
	if ((((66'sh3ffffffffffffffff >>> (8'sh32 <<< 4'shf)) & (W0131[6'h19] ? (66'sh1169fc5f7822a56b4 <<< 8'shff) : (~ 66'sh3ffffffffffffffff))) >>> (W0096 <<< W0040)) != 66'sh0) if (check) $stop;
	if ((~ $signed(W0132[125:3])) != 123'sh022cbf140000000021e199cf4e4f2fe) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (((((111'sh0 | 111'sh0) <<< W0096) | ((((111'sh0)==111'h0 ? 111'sh0:(111'sh0000000000010000000000000000 % 111'sh0)))==111'h0 ? 111'sh0:((111'sh7fffffffffffffffffffffffffff >>> 8'sh0) / ((111'sh0)==111'h0 ? 111'sh0:(111'sh0000000000010000000000000000 % 111'sh0))))) >>> ((8'sh0)==8'h0 ? 8'sh0:((W0015 <<< (4'shf & 4'sh5)) / 8'sh0))) != 111'sh0) if (check) $stop;
	if (58'sh000000021435d6c != 58'sh000000021435d6c) if (check) $stop;
   end
	//============================================================
   always @(check or W0015 or W0111 or W0040) begin : Block61
	W0133 = ((63'sh7fffffffffffffff & 63'sh7fffffffffffffff) >>> (1'h1 ? 7'sh0 : 7'sh0a));
	if (((((((~ 101'sh1fffffffffffffffffffffffff))==101'h0 ? 101'sh0:(((101'sh07801e45c800000000ffffffff)==101'h0 ? 101'sh0:(101'sh1fffffffffffffffffffffffff / 101'sh07801e45c800000000ffffffff)) / (~ 101'sh1fffffffffffffffffffffffff))) <<< (W0015 >>> W0040)))==101'h0 ? 101'sh0:(101'sh00000000000000000000000001 % ((((~ 101'sh1fffffffffffffffffffffffff))==101'h0 ? 101'sh0:(((101'sh07801e45c800000000ffffffff)==101'h0 ? 101'sh0:(101'sh1fffffffffffffffffffffffff / 101'sh07801e45c800000000ffffffff)) / (~ 101'sh1fffffffffffffffffffffffff))) <<< (W0015 >>> W0040)))) != 101'sh0) if (check) $stop;
	if ((W0133 >>> (((W0111)==7'h0 ? 7'sh0:((7'sh7f >>> 4'shd) % W0111)) >>> W0040)) != 63'sh7fffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(check or W0061) begin : Block62
	W0136 = (1'h1 ? 77'h0 : ((77'h0)==77'h0 ? 77'h0:(77'h1fffffffffffffffffff % 77'h0)));
	W0135 = 112'shffffffffffffffffffffffffffff;
	W0134 = W0135[111:72];
	if (((((({8{5'sh01}})==40'h0 ? 40'h0:((40'h0 & 40'h0bd1a118bf) % {8{5'sh01}})))==40'h0 ? 40'h0:(W0134 % (({8{5'sh01}})==40'h0 ? 40'h0:((40'h0 & 40'h0bd1a118bf) % {8{5'sh01}})))) & W0136[76:37]) != 40'h0) if (check) $stop;
	if (W0061 != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0139 <= 115'sh7ffffffffffffffffffffffffffff;
   end
   always @(posedge clk) begin
	W0138 <= W0139[114:1];
   end
   always @(posedge clk) begin
	W0137 <= (W0120 - W0138[113:113]);
   end
   always @(posedge clk) begin
	if (((((25'sh0 >>> 6'sh0) >>> (6'sh3f <<< 4'sh2)) >>> (W0090 <<< (4'sh7 >>> 3'sh7))) <= (((25'sh0 <<< 6'sh3f) >>> (6'sh0 >>> 4'shf)) >>> W0090)) != 1'h1) if (check) $stop;
	if (W0137 != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0143 <= ((128'sh0 >>> 8'sh01) >>> 8'sh01);
   end
   always @(posedge clk) begin
	W0142 <= W0143[126-:127];
   end
   always @(posedge clk) begin
	W0141 <= (~ 7'sh0);
   end
   always @(posedge clk) begin
	W0140 <= ((((42'sh3ff00000000)==42'h0 ? 42'sh0:(42'sh00000000001 / 42'sh3ff00000000)) <<< 7'sh7f) <<< W0141);
   end
   always @(posedge clk) begin
	if (W0140[41:40] != 2'h0) if (check) $stop;
	if (W0142[126:95] != 32'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0145 <= 91'sh0fc147500000000a1a6dc1c;
   end
   always @(posedge clk) begin
	W0144 <= W0145;
   end
   always @(posedge clk) begin
	if ($signed((W0144[90:90] ? 95'sh000000000000000000000001 : 95'sh0)) != 95'sh0) if (check) $stop;
	if (84'shfffffffffffffffffffff != 84'shfffffffffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(check or W0015) begin : Block66
	W0146 = 53'sh1fffffffffffff;
	if (((((98'sh3ffffffffffffffffffffffff)==98'h0 ? 98'sh0:((98'sh2fffffffffffffffff4e32117 >>> 8'sh45) % 98'sh3ffffffffffffffffffffffff)) >>> (($signed(8'hff))==8'h0 ? 8'sh0:(W0015 % $signed(8'hff)))) >>> 8'sh0) != 98'sh0) if (check) $stop;
	if ({1{(((W0146 | ((53'sh1fffffffffffff)==53'h0 ? 53'sh0:(53'sh0 / 53'sh1fffffffffffff))))==53'h0 ? 53'sh0:((($signed(53'h0ba454f928a5aa))==53'h0 ? 53'sh0:((~ 53'sh0) % $signed(53'h0ba454f928a5aa))) % (W0146 | ((53'sh1fffffffffffff)==53'h0 ? 53'sh0:(53'sh0 / 53'sh1fffffffffffff)))))}} != 53'h0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block67
	if ((((((18'sh3ffff <<< 6'sh01))==18'h0 ? 18'sh0:((18'sh0 >>> 6'sh01) % (18'sh3ffff <<< 6'sh01))) <<< (((6'sh01)==6'h0 ? 6'sh0:(6'sh3f / 6'sh01)) <<< 4'shc)) === (18'h0 << ((1'h0 ? 6'h01 : 6'h0) >> (~ 4'h2)))) != 1'h1) if (check) $stop;
	if (32'hda3f2a15 != 32'hda3f2a15) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0147 <= (76'shbc2ffffffff61887cef >>> W0096);
   end
   always @(posedge clk) begin
	if (57'sh1ded308896e764f != 57'sh1ded308896e764f) if (check) $stop;
	if ((W0147[75:41] << 7'h0) != 35'h5e17fffff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0149 <= (96'shffffffffffffffffffffffff + 96'shffffffffffffffffffffffff);
   end
   always @(posedge clk) begin
	W0148 <= (W0149 >>> (W0096 <<< W0105));
   end
   always @(posedge clk) begin
	if ($signed(W0053) != 2'sh0) if (check) $stop;
	if (W0148[95:17] != 79'h7fffffffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(check or W0053 or W0030 or W0002) begin : Block70
	W0150 = (- W0030);
	if (W0053 != 2'sh0) if (check) $stop;
	if (((64'hffffffffffffffff)==64'h0 ? 64'h0:(W0150[((1'h0 <  1'h0) ? W0002 : W0002)+:64] / 64'hffffffffffffffff)) != 64'h0) if (check) $stop;
   end
	//============================================================
   always @(check or W0120) begin : Block71
	W0151 = 6'sh0;
	if ((~ (31'sh00000001 >>> (W0151 >>> ((4'shf)==4'h0 ? 4'sh0:(4'sh0 % 4'shf))))) != 31'sh7ffffffe) if (check) $stop;
	if (W0120 != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block72
	W0155 = ((((35'sh7ffffffff <<< 7'sh01) & (35'sh7ffffffff | 35'sh0)))==35'h0 ? 35'sh0:(((((35'sh75f98c1bf)==35'h0 ? 35'sh0:(35'sh4233277ef / 35'sh75f98c1bf)))==35'h0 ? 35'sh0:(((35'sh6ffffffff)==35'h0 ? 35'sh0:(35'sh1e1da29e7 % 35'sh6ffffffff)) % ((35'sh75f98c1bf)==35'h0 ? 35'sh0:(35'sh4233277ef / 35'sh75f98c1bf)))) / ((35'sh7ffffffff <<< 7'sh01) & (35'sh7ffffffff | 35'sh0))));
	W0154 = 35'sh700000000;
	W0153 = W0154;
	W0152 = W0153[3+:32];
   end
   always @(posedge clk) begin : Block72Check
	if (((W0152[31:0])==32'h0 ? 32'h0:(32'h5d01711b / W0152[31:0])) != 32'h0) if (check) $stop;
	if (W0155[5'h0+:1] != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (W0137 != 1'h1) if (check) $stop;
	if (W0032 != 64'shfffffffe00000001) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0158 <= 108'sh000000000000000000000000001;
   end
   always @(posedge clk) begin
	W0157 <= W0158[107:1];
   end
   always @(posedge clk) begin
	W0156 <= ((121'sh1ffffffb6cbffd8ffffffff00000001)==121'h0 ? 121'sh0:(121'sh000000003d719e8ffffffffffffffff % 121'sh1ffffffb6cbffd8ffffffff00000001));
   end
   always @(posedge clk) begin
	if (W0037 != 31'sh7fffffff) if (check) $stop;
	if (({43'h0,(1'h1 ? W0133 : W0133)} & (W0156[120:15] >> W0157[40-:8])) != 106'h0000000000033d1ffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(check or W0003 or W0011) begin : Block75
	W0164 = W0003;
	W0163 = W0164[99-:87];
	W0162 = 117'sh1fffffffffffffffffffffffffffff;
	W0161 = ((96'hffffffffffffffffffffffff << 8'h01) + W0162[116:21]);
	W0160 = W0011;
	W0159 = ((60'sh000000000000001)==60'h0 ? 60'sh0:(60'sh000000000000001 / 60'sh000000000000001));
   end
   always @(posedge clk) begin : Block75Check
	if (((W0159[59:17] >> W0160) || 64'h000000000432c7fd) != 1'h1) if (check) $stop;
	if ((W0161 || W0163[3+:84]) != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(check or W0061) begin : Block76
	W0168 = (18'sh00001 - 18'sh3ffff);
	W0167 = (W0061 ? W0168 : (((18'sh0 & 18'sh17c61))==18'h0 ? 18'sh0:(18'sh0d0f6 / (18'sh0 & 18'sh17c61))));
	W0166 = (87'sh0 >>> 8'shff);
	W0165 = {W0166[86:63],((41'sh1ffffffffff)==41'h0 ? 41'sh0:((41'sh1ffffffffff <<< 7'sh1a) / 41'sh1ffffffffff))};
   end
   always @(posedge clk) begin : Block76Check
	if (W0165[64:64] != 1'h0) if (check) $stop;
	if (W0167[17:17] != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0171 <= (97'sh1ffffffffffffffffffffffff >>> (8'shff <<< 4'shf));
   end
   always @(posedge clk) begin
	W0170 <= (~ (118'sh0 >>> 8'sh01));
   end
   always @(posedge clk) begin
	W0169 <= (96'sh2eb5a3feffffffffa74f99bd - 96'sh00000001865cd906ffffffff);
   end
   always @(posedge clk) begin
	if ((((W0169)==96'h0 ? 96'sh0:((96'sh13b76419e266c572464d6815 ^ W0149) / W0169)) <<< W0015) != 96'sh0) if (check) $stop;
	if (((W0171[96:33])==64'h0 ? 64'h0:(W0170[117:54] % W0171[96:33])) != 64'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0174 <= 117'h1fffffffffffffffffffffffffffff;
   end
   always @(posedge clk) begin
	W0173 <= (((117'h000000000000000000000000000001)==117'h0 ? 117'h0:(117'h0 / 117'h000000000000000000000000000001)) & W0174);
   end
   always @(posedge clk) begin
	W0172 <= W0173[116:22];
   end
   always @(posedge clk) begin
	if (W0137 != 1'h1) if (check) $stop;
	if (W0172[6'h01] != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0178 <= 68'shf00000000ffffffff;
   end
   always @(posedge clk) begin
	W0177 <= W0178[67:30];
   end
   always @(posedge clk) begin
	W0176 <= W0177[37:37];
   end
   always @(posedge clk) begin
	W0175 <= (({23{1'h1}})==23'h0 ? 23'h0:((~ 23'h7fffff) / {23{1'h1}}));
   end
   always @(posedge clk) begin
	if ((~ (((((85'sh0 >>> 8'sh06))==85'h0 ? 85'sh0:(85'sh000000ffffffff0c94e8cc / (85'sh0 >>> 8'sh06))))==85'h0 ? 85'sh0:((- 85'sh18109300000000ffffffff) % (((85'sh0 >>> 8'sh06))==85'h0 ? 85'sh0:(85'sh000000ffffffff0c94e8cc / (85'sh0 >>> 8'sh06)))))) != 85'sh1fffffffffffffffffffff) if (check) $stop;
	if ((W0175[16-:1] >> W0176) != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0180 <= 8'shff;
   end
   always @(posedge clk) begin
	W0179 <= ((W0120 ? (68'sh0 <<< 8'sh01) : (68'sh0 >>> 8'shff)) >>> (((8'shff)==8'h0 ? 8'sh0:(8'shff % 8'shff)) & W0180));
   end
   always @(posedge clk) begin
	if (105'sh1ffffffffffffffffffffffffff != 105'sh1ffffffffffffffffffffffffff) if (check) $stop;
	if (W0179[67:8] != 60'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0185 <= 5'h01;
   end
   always @(posedge clk) begin
	W0184 <= 43'h7ffffffffff;
   end
   always @(posedge clk) begin
	W0183 <= 59'sh7ffffffffffffff;
   end
   always @(posedge clk) begin
	W0182 <= (~ 128'sh0);
   end
   always @(posedge clk) begin
	W0181 <= W0182[W0183[52-:6]+:35];
   end
   always @(posedge clk) begin
	if ((W0047 >>> W0015) != 96'shffffffffffffffffffffffff) if (check) $stop;
	if ((W0181[25-:1] ^ W0184[(W0185 ^ ((5'h1f)==5'h0 ? 5'h0:(5'h01 / 5'h1f)))+:1]) != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block82
	W0186 = (((120'h0 << (8'h0 | 8'h0)))==120'h0 ? 120'h0:(120'h000000ec84af558ee1d84a00000000 % (120'h0 << (8'h0 | 8'h0))));
	if (38'sh3fffffffff != 38'sh3fffffffff) if (check) $stop;
	if (W0186[119:13] != 107'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (W0168 != 18'sh00002) if (check) $stop;
	if ((($signed((((124'h9b9af1e694338baffffffffdbdf2475 << 8'hff))==124'h0 ? 124'h0:((1'h1 ? 124'hfffffffffffffffffffffffffffffff : 124'h9ecb5e63d0fd22700000000d6312ec0) % (124'h9b9af1e694338baffffffffdbdf2475 << 8'hff)))))==124'h0 ? 124'sh0:(((((124'sh0)==124'h0 ? 124'sh0:(124'sh0 / 124'sh0)) ^ ((124'sh000000000000000ffffffff00000001)==124'h0 ? 124'sh0:(124'sh0 / 124'sh000000000000000ffffffff00000001))) >>> W0180) / $signed((((124'h9b9af1e694338baffffffffdbdf2475 << 8'hff))==124'h0 ? 124'h0:((1'h1 ? 124'hfffffffffffffffffffffffffffffff : 124'h9ecb5e63d0fd22700000000d6312ec0) % (124'h9b9af1e694338baffffffffdbdf2475 << 8'hff)))))) != 124'sh0) if (check) $stop;
   end
	//============================================================
   always @(check or W0015) begin : Block84
	W0187 = (- ((121'sh0000000ffffffffffffffff00000000 | 121'sh00000000000000027ab4e109b3bd2b5) >>> W0015));
	if (W0187[120:49] != 72'hffffff800000000000) if (check) $stop;
	if (((109'sh0d0ad5a17d4e2105991700000000)==109'h0 ? 109'sh0:(109'sh0 / 109'sh0d0ad5a17d4e2105991700000000)) != 109'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (28'hfffffff != 28'hfffffff) if (check) $stop;
	if (W0032 != 64'shfffffffe00000001) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0192 <= (3'sh7 | 3'sh0);
   end
   always @(posedge clk) begin
	W0191 <= (~ 9'h1ff);
   end
   always @(posedge clk) begin
	W0190 <= 123'sh7ffffff079f4d86000000009983636f;
   end
   always @(posedge clk) begin
	W0189 <= W0190[122:18];
   end
   always @(posedge clk) begin
	W0188 <= (~ 128'shffffffffffffffffffffffffffffffff);
   end
   always @(posedge clk) begin
	if ((W0188[113-:80] << (W0189[104:97] << W0191[8:5])) != 80'h0) if (check) $stop;
	if ((~ W0192[0-:1]) != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(check or W0054) begin : Block87
	W0193 = (((31'sh7fffffff >  31'h7fffffff) ? W0054 : W0054) - W0054);
	if (((28'shbf65019)==28'h0 ? 28'sh0:(28'sh0 / 28'shbf65019)) != 28'sh0) if (check) $stop;
	if (W0193 != 2'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0195 <= (31'sh00000001 >>> W0084);
   end
   always @(posedge clk) begin
	W0194 <= 35'sh600000000;
   end
   always @(posedge clk) begin
	if (W0194[6-:1] != 1'h0) if (check) $stop;
	if (W0195 != 31'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0196 <= W0176;
   end
   always @(posedge clk) begin
	if (W0196 != 1'h1) if (check) $stop;
	if (W0032 != 64'shfffffffe00000001) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (31'sh7fffffff != 31'sh7fffffff) if (check) $stop;
	if (((~ W0133) | ((W0133)==63'h0 ? 63'sh0:(((W0133)==63'h0 ? 63'sh0:((63'sh0000000000000001 <<< 7'sh53) % W0133)) % W0133))) != 63'sh0) if (check) $stop;
   end
	//============================================================
   always @(check or W0196 or W0002 or W0042) begin : Block91
	W0198 = 15'h0;
	W0197 = 111'sh0;
	if ((((W0196 << W0196))==1'h0 ? 1'h0:(1'h0 % (W0196 << W0196))) != 1'h0) if (check) $stop;
	if ((({{22{W0198[3'h7]}},(((64'shffffffffffffffff)==64'h0 ? 64'sh0:(64'sh2aafe03affffffff / 64'shffffffffffffffff)) >>> W0042)})==86'h0 ? 86'h0:(W0197[W0002+:86] % {{22{W0198[3'h7]}},(((64'shffffffffffffffff)==64'h0 ? 64'sh0:(64'sh2aafe03affffffff / 64'shffffffffffffffff)) >>> W0042)})) != 86'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0199 <= 25'sh1930f53;
   end
   always @(posedge clk) begin
	if ((((W0199)==25'h0 ? 25'sh0:(((95'h1792207dffffffff00000000 !== 95'sh7fffffffffffffffffffffff) ? ((25'sh0000001)==25'h0 ? 25'sh0:(25'sh0 / 25'sh0000001)) : (1'h1 ? 25'sh1ffffff : 25'sh0)) % W0199)) <<< W0151) != 25'sh0) if (check) $stop;
	if (75'h45708c934aad6da79b4 != 75'h45708c934aad6da79b4) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0201 <= 62'sh3fffffffffffffff;
   end
   always @(posedge clk) begin
	W0200 <= (1'h0 << 1'h1);
   end
   always @(posedge clk) begin
	if ((((W0200)==1'h0 ? 1'h0:(1'h1 / W0200)) ? ((62'sh3fffffffffffffff)==62'h0 ? 62'sh0:((W0201 >>> W0042) % 62'sh3fffffffffffffff)) : 62'sh0000000100000000) != 62'sh0000000100000000) if (check) $stop;
	if ((W0037 >>> W0084) != 31'sh7fffffff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0207 <= ((125'sh0 >>> (8'sh94 <<< 4'sh1)) - ((~ 125'sh0) >>> (8'sh0 >>> 4'sh6)));
   end
   always @(posedge clk) begin
	W0206 <= 99'sh0;
   end
   always @(posedge clk) begin
	W0205 <= W0206[79-:4];
   end
   always @(posedge clk) begin
	W0204 <= 29'h1f3fc1c3;
   end
   always @(posedge clk) begin
	W0203 <= {28'shf662aa6,55'sh12a8ed00000000};
   end
   always @(posedge clk) begin
	W0202 <= (($signed(128'hffffffffffffffffffffffffffffffff))==128'h0 ? 128'sh0:((128'shffffffffffffffffffffffffffffffff >>> 8'shff) % $signed(128'hffffffffffffffffffffffffffffffff)));
   end
   always @(posedge clk) begin
	if ((W0202[((((4'h0)==4'h0 ? 4'h0:(4'hf / 4'h0)))==4'h0 ? 4'h0:(((4'h0)==4'h0 ? 4'h0:(4'h1 % 4'h0)) % ((4'h0)==4'h0 ? 4'h0:(4'hf / 4'h0))))+:109] >> (W0203[W0204[28:23]+:8] << W0205)) != 109'h0) if (check) $stop;
	if (W0207 != 125'sh00000000000000000000000000000001) if (check) $stop;
   end
	//============================================================
   always @(check or W0151 or W0036 or W0017 or W0105) begin : Block95
	W0208 = (((105'sh000ffffffffffffffff50906cd4 <<< 8'sh0))==105'h0 ? 105'sh0:(((105'sh1ff84dad3b87c263736062a0982)==105'h0 ? 105'sh0:(105'sh1ffffffffff74d9a69a78dbe00c / 105'sh1ff84dad3b87c263736062a0982)) / (105'sh000ffffffffffffffff50906cd4 <<< 8'sh0)));
	if ((W0017 <<< (((W0151)==6'h0 ? 6'sh0:(6'sh01 % W0151)) >>> W0105)) != 32'shffffffff) if (check) $stop;
	if (((W0036)==95'h0 ? 95'h0:(W0208[104:10] % W0036)) != 95'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0209 <= (((101'sh0)==101'h0 ? 101'sh0:(101'sh0 / 101'sh0)) - 101'sh0000000000ffffffffffffffff);
   end
   always @(posedge clk) begin
	if (((~ (W0196 << 1'h1)) ? 101'sh008767606855af5f46ffffffff : W0209) != 101'sh008767606855af5f46ffffffff) if (check) $stop;
	if (W0083 != 32'sh0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block97
   end
   always @(posedge clk) begin : Block97Check
	if (32'sh0 != 32'sh0) if (check) $stop;
	if (96'shffffffffffffffffffffffff != 96'shffffffffffffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(check or W0196) begin : Block98
	W0211 = ((~ 1'h0) ? (111'sh0 >>> 8'sh0) : (111'sh0000ef79dda4ffffffffffffffff >>> 8'shff));
	W0210 = W0211[110:109];
   end
   always @(posedge clk) begin : Block98Check
	if (W0196 != 1'h1) if (check) $stop;
	if (W0210 != 2'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0216 <= 15'h0;
   end
   always @(posedge clk) begin
	W0215 <= W0216[9-:6];
   end
   always @(posedge clk) begin
	W0214 <= W0209;
   end
   always @(posedge clk) begin
	W0213 <= 98'sh0000000000000000000000001;
   end
   always @(posedge clk) begin
	W0212 <= {63{W0214[100:100]}};
   end
   always @(posedge clk) begin
	if (W0212[(W0213[97:93] << 4'h0)+:1] != 1'h1) if (check) $stop;
	if ((((~ W0215[5:5]))==1'h0 ? 1'h0:((W0037 == W0037) % (~ W0215[5:5]))) != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0219 <= 103'sh00000000000000000000000001;
   end
   always @(posedge clk) begin
	W0218 <= 103'sh0085bac6fde88fbe57a202d84c;
   end
   always @(posedge clk) begin
	W0217 <= ((((W0219)==103'h0 ? 103'sh0:((103'sh0 >>> 8'shff) % W0219)))==103'h0 ? 103'sh0:(((1'h1 | 1'h1) ? W0218 : (103'sh0 <<< 8'sh01)) / ((W0219)==103'h0 ? 103'sh0:((103'sh0 >>> 8'shff) % W0219))));
   end
   always @(posedge clk) begin
	if (W0133 != 63'sh7fffffffffffffff) if (check) $stop;
	if (W0217[102:102] != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0223 <= {3'h1,122'sh0};
   end
   always @(posedge clk) begin
	W0222 <= ((((99'sh7ffffffff00000000ffffffff)==99'h0 ? 99'sh0:(99'sh1ffffffffb5bae196a0f8ef2e % 99'sh7ffffffff00000000ffffffff)))==99'h0 ? 99'sh0:((1'h1 ? 99'sh0 : 99'sh0000000000000000000000001) % ((99'sh7ffffffff00000000ffffffff)==99'h0 ? 99'sh0:(99'sh1ffffffffb5bae196a0f8ef2e % 99'sh7ffffffff00000000ffffffff))));
   end
   always @(posedge clk) begin
	W0221 <= 105'sh18b7e03b2359874995a00000000;
   end
   always @(posedge clk) begin
	W0220 <= (~ 35'sh700000001);
   end
   always @(posedge clk) begin
	if ((W0220[(W0221[104:104] ? W0185 : ((5'h1f)==5'h0 ? 5'h0:(5'h0 % 5'h1f)))+:1] >> W0222[28-:1]) != 1'h1) if (check) $stop;
	if (W0223[124:61] != 64'h2000000000000000) if (check) $stop;
   end
	//============================================================
   always @(check or W0200) begin : Block102
	W0225 = (1'h0 ? 103'sh7f0000000000000000a932571f : 103'sh7fffffffffffffffffffffffff);
	W0224 = W0225[99-:99];
	if (((W0224[94-:95])==95'h0 ? 95'h0:(95'h7fffffffffffffffffffffff / W0224[94-:95])) != 95'h000000000000000000000001) if (check) $stop;
	if (W0200 != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(check or W0160) begin : Block103
   end
   always @(posedge clk) begin : Block103Check
	if ((((~ 119'sh7fffffffffffffffffffffffffffff) | (~ ((119'sh558215000000000000000000000001)==119'h0 ? 119'sh0:(119'sh6160ec5908bbfcffffffff19180b72 / 119'sh558215000000000000000000000001)))) & 119'sh0) != 119'sh0) if (check) $stop;
	if ((64'hffffffffffffffff << W0160) != 64'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (15'sh39b6 != 15'sh39b6) if (check) $stop;
	if (W0133 != 63'sh7fffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0228 <= 5'sh10;
   end
   always @(posedge clk) begin
	W0227 <= 5'sh1f;
   end
   always @(posedge clk) begin
	W0226 <= 5'sh0;
   end
   always @(posedge clk) begin
	if (52'sh0 != 52'sh0) if (check) $stop;
	if (((((W0227 <<< (4'shf >>> 3'sh1)) | (- W0228)))==5'h0 ? 5'sh0:(((W0226 >>> W0040) >>> W0105) / ((W0227 <<< (4'shf >>> 3'sh1)) | (- W0228)))) != 5'sh0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block106
	W0230 = (& (14'sh0001 >>> 5'sh1f));
	W0229 = 3'sh3;
	if ((W0229[(1'h0 ? {1{1'h0}} : (1'h1 | 1'h1))] << ({6'h0,4'sh1} !== 10'sh0)) != 1'h0) if (check) $stop;
	if ({1{W0230}} != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block107
	W0232 = 95'h0;
	W0231 = 128'h0;
	if (W0231 != 128'h0) if (check) $stop;
	if (((W0232[94:63])==32'h0 ? 32'h0:(32'hffffffff / W0232[94:63])) != 32'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0233 <= ((((14'sh3fff)==14'h0 ? 14'sh0:(14'sh0 % 14'sh3fff)))==14'h0 ? 14'sh0:(14'sh0 % ((14'sh3fff)==14'h0 ? 14'sh0:(14'sh0 % 14'sh3fff))));
   end
   always @(posedge clk) begin
	if (32'sh0 != 32'sh0) if (check) $stop;
	if ((14'sh3fff | W0233) != 14'sh3fff) if (check) $stop;
   end
	//============================================================
   always @(check or W0180) begin : Block109
	W0235 = W0180;
	W0234 = ($signed(((127'sh000000010000000065c23b2a00000001)==127'h0 ? 127'sh0:(127'sh00000000000000018a995eff00000000 / 127'sh000000010000000065c23b2a00000001))) >>> W0235);
   end
   always @(posedge clk) begin : Block109Check
	if (($signed(96'hffffffffffffffffffffffff) >>> W0180) != 96'shffffffffffffffffffffffff) if (check) $stop;
	if (W0234[126:126] != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block110
	W0236 = 37'sh1fffffffff;
   end
   always @(posedge clk) begin : Block110Check
	if (((((((W0236)==37'h0 ? 37'sh0:((37'sh137942ceb2 <<< 7'sh01) % W0236)))==37'h0 ? 37'sh0:(37'sh0 / ((W0236)==37'h0 ? 37'sh0:((37'sh137942ceb2 <<< 7'sh01) % W0236)))))==37'h0 ? 37'sh0:(37'sh1fffffffff / ((((W0236)==37'h0 ? 37'sh0:((37'sh137942ceb2 <<< 7'sh01) % W0236)))==37'h0 ? 37'sh0:(37'sh0 / ((W0236)==37'h0 ? 37'sh0:((37'sh137942ceb2 <<< 7'sh01) % W0236)))))) != 37'sh0) if (check) $stop;
	if ((47'sh627035bf7a97 & ((((47'sh7fff00000000 >>> 7'sh7f) >>> (7'sh7f | 7'sh0)))==47'h0 ? 47'sh0:(47'sh7fffffffffff / ((47'sh7fff00000000 >>> 7'sh7f) >>> (7'sh7f | 7'sh0))))) != 47'sh000000000001) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0239 <= 123'sh53fb225d8fa2187ffffffffffffffff;
   end
   always @(posedge clk) begin
	W0238 <= (119'sh000000ffffffff0000000000000000 ^ 119'sh7fffffffffffffffffffffffffffff);
   end
   always @(posedge clk) begin
	W0237 <= W0238[68-:1];
   end
   always @(posedge clk) begin
	if ((W0237 ? 21'sh000001 : (~ $signed(21'sh000001))) != 21'sh1ffffe) if (check) $stop;
	if ((~ W0239[122:60]) != 63'h2c04dda2705de780) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (W0031 != 64'shfffffffe00000001) if (check) $stop;
	if (((~| ((110'h0 >> 8'h0) != (110'sh00000000000000000000ffffffff >>> 8'shff))) << 1'h0) != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0242 <= 6'sh3f;
   end
   always @(posedge clk) begin
	W0241 <= 67'sh7ffffffffee0efff1;
   end
   always @(posedge clk) begin
	W0240 <= 50'sh0;
   end
   always @(posedge clk) begin
	if ((((50'sh0000078a01e1c)==50'h0 ? 50'sh0:((W0240 >>> ((7'sh7f)==7'h0 ? 7'sh0:(7'sh01 % 7'sh7f))) % 50'sh0000078a01e1c)) ^ (((50'sh2b919ca68fa68 | ((50'sh0)==50'h0 ? 50'sh0:(50'sh0000000000001 / 50'sh0))))==50'h0 ? 50'sh0:((W0241[66:66] ? ((50'sh0)==50'h0 ? 50'sh0:(50'sh00000ffffffff / 50'sh0)) : ((50'sh0)==50'h0 ? 50'sh0:(50'sh0 / 50'sh0))) / (50'sh2b919ca68fa68 | ((50'sh0)==50'h0 ? 50'sh0:(50'sh0000000000001 / 50'sh0)))))) != 50'sh0) if (check) $stop;
	if (((((26'sh3ffffff <<< 6'sh01) >>> W0242) <<< (W0151 | W0090)) <<< 6'sh0) != 26'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0243 <= (W0061 ? (1'h1 ? 32'hffffffff : 32'h2c0ee208) : ((32'h0)==32'h0 ? 32'h0:(32'h0 % 32'h0)));
   end
   always @(posedge clk) begin
	if (W0031 != 64'shfffffffe00000001) if (check) $stop;
	if ((W0243 << 6'h3f) != 32'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0247 <= ((75'sh0)==75'h0 ? 75'sh0:(75'sh0 % 75'sh0));
   end
   always @(posedge clk) begin
	W0246 <= 3'sh7;
   end
   always @(posedge clk) begin
	W0245 <= 4'shf;
   end
   always @(posedge clk) begin
	W0244 <= (8'sh0 - 8'sh8d);
   end
   always @(posedge clk) begin
	if ((((- (1'h0 ? 109'sh00005cd67561a89d641e00000001 : 109'sh0000000000000000000000000001)) <<< W0235) >>> (W0244 >>> (W0245 <<< W0246))) != 109'sh0) if (check) $stop;
	if ((82'sh3ffffffffffffffffffff <<< (W0247[(6'h0 >> 4'h0)+:1] ? (((8'shff)==8'h0 ? 8'sh0:(8'sh5b % 8'shff)) >>> (~ 4'sh0)) : ((W0015)==8'h0 ? 8'sh0:((8'sh01 >>> 4'shf) / W0015)))) != 82'sh3ffffffffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(check or W0237) begin : Block116
	if (W0237 != 1'h0) if (check) $stop;
	if (57'sh0 != 57'sh0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block117
	if ({8'h0,((56'sh00000000000001)==56'h0 ? 56'sh0:(((56'sh00000000000001 >>> 7'sh7f) <<< (7'sh3f >>> 4'sh0)) / 56'sh00000000000001))} != 64'h0) if (check) $stop;
	if (63'sh0 != 63'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (W0052 != 2'sh0) if (check) $stop;
	if (((96'shffffffffffffffffffffffff)==96'h0 ? 96'sh0:(W0047 % 96'shffffffffffffffffffffffff)) != 96'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0252 <= 96'h0;
   end
   always @(posedge clk) begin
	W0251 <= W0252[95:41];
   end
   always @(posedge clk) begin
	W0250 <= 93'sh0;
   end
   always @(posedge clk) begin
	W0249 <= 43'h7ffffffffff;
   end
   always @(posedge clk) begin
	W0248 <= (((28'shfffffff <<< 6'sh3f) >>> (- 6'sh1c)) * (- (28'shfffffff >>> 6'sh0)));
   end
   always @(posedge clk) begin
	if (W0248 != 28'sh0) if (check) $stop;
	if ((W0249[42:29] & ((((1'h0 ? 14'h3fff : 14'h0))==14'h0 ? 14'h0:(W0250[92:79] % (1'h0 ? 14'h3fff : 14'h0))) >> W0251[54:50])) != 14'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0254 <= 79'sh7fff87182181ffffffff;
   end
   always @(posedge clk) begin
	W0253 <= W0028;
   end
   always @(posedge clk) begin
	if (W0253[W0254[78:74]] != 1'h0) if (check) $stop;
	if ((W0195 >>> W0151) != 31'sh0) if (check) $stop;
   end
	//============================================================
   always @(check or W0137) begin : Block121
	W0255 = (((~ (127'h0 << 8'hd7)))==127'h0 ? 127'h0:(127'h0 % (~ (127'h0 << 8'hd7))));
	if (W0255[126:0] != 127'h0) if (check) $stop;
	if (W0137 != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0259 <= ((81'sh1ffffffffffffffffffff >>> 8'shff) >>> ((8'shff)==8'h0 ? 8'sh0:(8'sh01 / 8'shff)));
   end
   always @(posedge clk) begin
	W0258 <= ((~ 113'h1ffffffffffffffffffffffffffff) >> W0125);
   end
   always @(posedge clk) begin
	W0257 <= W0196;
   end
   always @(posedge clk) begin
	W0256 <= (78'sh0001000000014a8f216b <<< 8'sh01);
   end
   always @(posedge clk) begin
	if ($unsigned($signed(W0256)) != 78'h000200000002951e42d6) if (check) $stop;
	if ((W0257 ? W0258[112:49] : W0259[80:17]) != 64'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0260 <= $unsigned((((36'sh9627e9d6a)==36'h0 ? 36'sh0:(36'sh0a9f0c0a5 / 36'sh9627e9d6a)) & (1'h1 ? 36'sh0 : 36'sh6ffffffff)));
   end
   always @(posedge clk) begin
	if (W0133 != 63'sh7fffffffffffffff) if (check) $stop;
	if (W0260[35:21] != 15'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0262 <= (114'sh0 >>> 8'shff);
   end
   always @(posedge clk) begin
	W0261 <= W0262[113:11];
   end
   always @(posedge clk) begin
	if ($signed(W0261[102:71]) != 32'sh0) if (check) $stop;
	if (20'sh0 != 20'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0266 <= 31'sh7fffffff;
   end
   always @(posedge clk) begin
	W0265 <= 35'sh0;
   end
   always @(posedge clk) begin
	W0264 <= ((128'sh62aa887fd0add0ee000000009f6f690b)==128'h0 ? 128'sh0:(128'sh00000000000000000000000000000001 / 128'sh62aa887fd0add0ee000000009f6f690b));
   end
   always @(posedge clk) begin
	W0263 <= (W0264[59-:48] * (((48'hffffffffffff >> 7'h77))==48'h0 ? 48'h0:((~ 48'h0) % (48'hffffffffffff >> 7'h77))));
   end
   always @(posedge clk) begin
	if (W0263 != 48'h0) if (check) $stop;
	if ((~ W0265[W0266[11-:5]+:1]) != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(check or W0243 or W0242) begin : Block126
	W0269 = (128'shffffffffffffffffffffffffffffffff >>> 8'sh0);
	W0268 = (1'h1 ? 51'sh00000e748356c : 51'sh7ffff00000000);
	W0267 = {W0268[(4'h9 | 4'h0)+:23],W0269[5'h01+:68]};
   end
   always @(posedge clk) begin : Block126Check
	if ((W0243 >> $unsigned((~ W0242))) != 32'hffffffff) if (check) $stop;
	if (W0267[17-:1] != 1'h1) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0270 <= (((((19'sh7ffff >>> 6'sh3f))==19'h0 ? 19'sh0:(((19'sh0)==19'h0 ? 19'sh0:(19'sh00001 / 19'sh0)) / (19'sh7ffff >>> 6'sh3f))))==19'h0 ? 19'sh0:(19'sh0 / (((19'sh7ffff >>> 6'sh3f))==19'h0 ? 19'sh0:(((19'sh0)==19'h0 ? 19'sh0:(19'sh00001 / 19'sh0)) / (19'sh7ffff >>> 6'sh3f)))));
   end
   always @(posedge clk) begin
	if ($signed(W0161) != 96'shfffffffffffffffffffffffd) if (check) $stop;
	if (W0270[17-:18] != 18'h0) if (check) $stop;
   end
	//============================================================
   always @(check or W0196 or W0219) begin : Block128
	W0277 = 6'h3f;
	W0276 = W0219;
	W0275 = (((67'sh7ffffffffffffffff >>> 8'shff))==67'h0 ? 67'sh0:(67'sh7ffffffffffffffff % (67'sh7ffffffffffffffff >>> 8'shff)));
	W0274 = (((17'h0)==17'h0 ? 17'h0:(17'h0 / 17'h0)) * 17'h1ffff);
	W0273 = 35'h000000001;
	W0272 = 83'h51274ffffffffffffffff;
	W0271 = 54'sh00000000000001;
   end
   always @(posedge clk) begin : Block128Check
	if (((W0274)==17'h0 ? 17'h0:((((W0273[5'h01] ? (17'h0 >> 6'h24) : (17'h00001 >> 6'h30)))==17'h0 ? 17'h0:(((W0272[6'h3f+:17])==17'h0 ? 17'h0:(W0271[53:37] / W0272[6'h3f+:17])) % (W0273[5'h01] ? (17'h0 >> 6'h24) : (17'h00001 >> 6'h30)))) / W0274)) != 17'h0) if (check) $stop;
	if ((W0275[W0276[W0277+:6]+:1] << W0196) != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0280 <= W0120;
   end
   always @(posedge clk) begin
	W0279 <= (123'sh000000096e9e0b0ffffffff00000000 | 123'sh0000000fec7862400000000c7107e4a);
   end
   always @(posedge clk) begin
	W0278 <= (W0279[(6'h0 << 4'hf)+:1] ? ((1'h1 ? 10'sh3ff : 10'sh0) <<< W0228) : 10'sh3ff);
   end
   always @(posedge clk) begin
	if (W0278[9:9] != 1'h1) if (check) $stop;
	if (W0280[0:0] != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0282 <= {28'h0,22'h0};
   end
   always @(posedge clk) begin
	W0281 <= W0282;
   end
   always @(posedge clk) begin
	if (((1'h1)==1'h0 ? 1'h0:(W0281[49:49] % 1'h1)) != 1'h0) if (check) $stop;
	if ((- (~ 73'sh1ff0000000100000000)) != 73'sh1ff0000000100000001) if (check) $stop;
   end
	//============================================================
   always @(check or W0244 or W0015) begin : Block131
	if (95'h0 != 95'h0) if (check) $stop;
	if (((- ((1'h0 ? 69'sh1f000000005f6fd955 : 69'sh0) <<< W0015)) & (((69'sh1fffffffff6a435651 >>> W0244))==69'h0 ? 69'sh0:(((69'sh1fffffffffffffffff >>> 8'sh01) >>> (8'sh01 >>> 4'sh0)) % (69'sh1fffffffff6a435651 >>> W0244)))) != 69'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0285 <= 95'h7fffffffffffffffffffffff;
   end
   always @(posedge clk) begin
	W0284 <= {W0285,(33'h0ffffffff & 33'h1101dee12)};
   end
   always @(posedge clk) begin
	W0283 <= W0284[(- 5'h06)+:79];
   end
   always @(posedge clk) begin
	if (W0283[W0277] != 1'h1) if (check) $stop;
	if (54'sh00000000000001 != 54'sh00000000000001) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0288 <= 2'sh3;
   end
   always @(posedge clk) begin
	W0287 <= 1'h0;
   end
   always @(posedge clk) begin
	W0286 <= W0109;
   end
   always @(posedge clk) begin
	if ({41{W0286[20-:1]}} != 41'h0) if (check) $stop;
	if (((((19'sh43ea7)==19'h0 ? 19'sh0:((19'sh0 >>> 6'sh0) % 19'sh43ea7)) && (W0287 ? ((64'sh0)==64'h0 ? 64'sh0:(64'sh2117d19387012c11 % 64'sh0)) : (64'sh0 >>> 7'sh6b))) ? W0288 : W0054) != 2'sh0) if (check) $stop;
   end
	//============================================================
   always @(check or W0207 or W0099) begin : Block134
	W0289 = (((W0207 >>> (8'sh0 | 8'she4)))==125'h0 ? 125'sh0:(125'sh1fffffff000000012f126cb600000000 % (W0207 >>> (8'sh0 | 8'she4))));
	if (W0099 != 20'sh0) if (check) $stop;
	if (W0289[124:34] != 91'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if ((((((- 31'sh00000001) >>> 6'sh0))==31'h0 ? 31'sh0:((((31'sh7fffffff | 31'sh7fffffff))==31'h0 ? 31'sh0:((31'sh00000001 >>> 6'sh12) / (31'sh7fffffff | 31'sh7fffffff))) / ((- 31'sh00000001) >>> 6'sh0))) >>> W0090) != 31'sh0) if (check) $stop;
	if (52'shfffff00000000 != 52'shfffff00000000) if (check) $stop;
   end
	//============================================================
   always @(check or W0104 or W0015) begin : Block136
	W0296 = $unsigned(W0104);
	W0295 = (128'sh0000000100000000d0ed7551a8e8b0f8 >>> W0015);
	W0294 = 128'sh0000000000000000fffffffffe02e239;
	W0293 = W0294[2'h3+:121];
	W0292 = 121'sh1906da100000001ffffffff00000000;
	W0291 = W0292;
	W0290 = ((W0293[120:8])==113'h0 ? 113'h0:(W0291[120:8] % W0293[120:8]));
	if (W0290[112:112] != 1'h0) if (check) $stop;
	if ((W0295[122-:121] ^ W0296[121:1]) != 121'h1ffffffbfffffffcbc4a2ab95c5d3c1) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0303 <= 7'sh7f;
   end
   always @(posedge clk) begin
	W0302 <= W0168;
   end
   always @(posedge clk) begin
	W0301 <= (~ 27'sh0);
   end
   always @(posedge clk) begin
	W0300 <= ((((55'sh655f9bffffffff)==55'h0 ? 55'sh0:(55'sh7fffff7d8969a5 / 55'sh655f9bffffffff)) <<< W0303) <<< W0141);
   end
   always @(posedge clk) begin
	W0299 <= ((111'sh7fff000000010000000065b2bace ^ 111'sh0) >>> (8'shba <<< 4'sh0));
   end
   always @(posedge clk) begin
	W0298 <= 79'sh7fffffffffffffffffff;
   end
   always @(posedge clk) begin
	W0297 <= W0298[78:20];
   end
   always @(posedge clk) begin
	if (((W0196 ? ((((59'h7ffffffffffffff)==59'h0 ? 59'h0:(59'h0 % 59'h7ffffffffffffff)))==59'h0 ? 59'h0:((59'h0 << 7'h01) / ((59'h7ffffffffffffff)==59'h0 ? 59'h0:(59'h0 % 59'h7ffffffffffffff)))) : W0297) | W0299[(- (5'h0 >> 4'h1))+:59]) != 59'h7ffffffffffffff) if (check) $stop;
	if (W0300[((W0302[17:14])==4'h0 ? 4'h0:(W0301[26:23] / W0302[17:14]))+:32] != 32'h0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0304 <= (($unsigned((111'h7fffffffffffffffffffffffffff | 111'h7fffffffffffffffffffffffffff)))==111'h0 ? 111'h0:(111'h7fffffffffffffffffffffffffff % $unsigned((111'h7fffffffffffffffffffffffffff | 111'h7fffffffffffffffffffffffffff))));
   end
   always @(posedge clk) begin
	if (W0304[110:7] != 104'h0) if (check) $stop;
	if (W0037 != 31'sh7fffffff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if ((((W0133 <<< ((W0111)==7'h0 ? 7'sh0:((7'sh01 ^ 7'sh7f) / W0111))))==63'h0 ? 63'sh0:((W0133 >>> (W0111 <<< (4'sh0 | 4'shf))) % (W0133 <<< ((W0111)==7'h0 ? 7'sh0:((7'sh01 ^ 7'sh7f) / W0111))))) != 63'sh0) if (check) $stop;
	if ($unsigned((((21'sh0 | 21'sh000001) <<< W0090) <<< 6'sh3f)) != 21'h0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block140
	W0306 = 116'sh000004a144132ffffffffffffffff;
	W0305 = (((W0306[115:19])==97'h0 ? 97'h0:(97'h1ffffffffffffffffffffffff / W0306[115:19])) ^ {66'h0,31'sh0});
	if (W0305[96:54] != 43'h0) if (check) $stop;
	if (69'sh000000000000000001 != 69'sh000000000000000001) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (((W0032)==64'h0 ? 64'sh0:(64'sh7e2aefddd3bac6f5 / W0032)) != 64'shffffffffc0ea8811) if (check) $stop;
	if ((W0109 >>> 8'sh0) != 67'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (32'shffffffff != 32'shffffffff) if (check) $stop;
	if (2'sh0 != 2'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	W0308 <= 23'sh283d11;
   end
   always @(posedge clk) begin
	W0307 <= (W0308[4'h0] ? (20'h0 << 6'h0) : {15'h0,5'h0});
   end
   always @(posedge clk) begin
	if (W0120 != 1'h0) if (check) $stop;
	if ((W0307[19:19] && (W0195 >>> W0084)) != 1'h0) if (check) $stop;
   end
	//============================================================
   always @(check or W0003) begin : Block144
	W0311 = W0003;
	W0310 = W0311;
	W0309 = 86'h0;
	if (W0309 != 86'h0) if (check) $stop;
	if (W0310[2+:126] != 126'h3fffffffffffffffffffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block145
	if (63'sh0 != 63'sh0) if (check) $stop;
	if (100'sh0 != 100'sh0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block146
	W0312 = (1'h1 ? {52'h0,(2'sh3 <<< 2'sh3)} : ((54'h3fffff5dd55547 << 7'h7f) << 7'h0));
	if (97'sh1ffffffffd48a45d68db4e037 != 97'sh1ffffffffd48a45d68db4e037) if (check) $stop;
	if (W0312 != 54'h0) if (check) $stop;
   end
	//============================================================
   always @(check) begin : Block147
	W0315 = (111'sh0 * 111'sh0);
	W0314 = ((111'sh4ee300000000ffffffff00000000)==111'h0 ? 111'sh0:(111'sh0 / 111'sh4ee300000000ffffffff00000000));
	W0313 = (W0314 + W0315);
	if ((~ 95'h7fffffffffffffffffffffff) != 95'h0) if (check) $stop;
	if (W0313 != 111'sh0) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (((W0169)==96'h0 ? 96'sh0:(W0149 / W0169)) != 96'sh0) if (check) $stop;
	if (64'shffffffffffffffff != 64'shffffffffffffffff) if (check) $stop;
   end
	//============================================================
   always @(posedge clk) begin
	if (1'h0 != 1'h0) if (check) $stop;
	if (((W0292 >>> ((8'sh82)==8'h0 ? 8'sh0:(W0180 / 8'sh82))) <<< ((((8'shff <<< 4'sh1))==8'h0 ? 8'sh0:(W0096 / (8'shff <<< 4'sh1))) >>> ((W0105)==4'h0 ? 4'sh0:(4'sh0 % W0105)))) != 121'sh1906da100000001ffffffff00000000) if (check) $stop;
   end
	//============================================================
   always @(check or W0003) begin : Block150
	W0318 = (81'sh00000000000009787cfbe - 81'sh1ffff900819b062834600);
	W0317 = (W0318 - 81'sh0cabb9992e90800000000);
	W0316 = W0003;
	if (W0316[123-:124] != 124'hfffffffffffffffffffffffffffffff) if (check) $stop;
	if (W0317 != 81'sh13544d664fd48350489be) if (check) $stop;
   end

   reg done; initial done=1'b0;
   reg ddone; initial ddone=1'b0;
   always @(posedge clk) begin
      if (check) begin
         done <= 1'b1;
      end
      if (done && !ddone) begin
         ddone <= 1'b1;
         $write("*-* All Finished *-*\n");
      end
   end

   parameter [31:0] CYCLES /*verilator public*/ = 205;
endmodule
